`define DLY #1
//`define SIMULATION
`ifndef SIMULATION
  `define TEST_PAT0
//`define TEST_PAT1
//`define TEST_PAT2
//`define TEST_PAT3
`endif

module pic_gen(
    // global signals
    clk                 , // <i>  1b, global clock
    rstn                , // <i>  1b, global reset, active low
    // picture data output
    pic_hsync           , // <o>  1b, picture hsync
    pic_vsync           , // <o>  1b, picture vsync
    pic_dat_en          , // <o>  1b, picture data enable
    pic_data              // <o> 24b, picture data
    );

  // global signals
  input         clk                 ; // <i>  1b, global clock
  input         rstn                ; // <i>  1b, global reset, active low
  // picture data output
  output        pic_hsync           ; // <o>  1b, picture hsync
  output        pic_vsync           ; // <o>  1b, picture vsync
  output        pic_dat_en          ; // <o>  1b, picture data enable
  output [23:0] pic_data            ; // <o> 24b, picture data

  reg   [3:0]   clk_div             ;

  reg   [10:0]  hcnt                ;
  reg   [10:0]  vcnt                ;

`ifndef SIMULATION
  reg   [23:0]  pic_data            ;
`endif

`ifdef TEST_PAT0
  wire  [5:0]   pic_addr            ;
`elsif TEST_PAT1
  wire  [12:0]  pic_addr            ;
`elsif TEST_PAT2
`elsif TEST_PAT3
`endif

`ifdef SIMULATION
  reg   [23:0]  bmp_data_mem[0:2073599];
`endif

`ifdef SIMULATION
  parameter HTOTAL  = 2048;
  parameter VTOTAL  = 1400;
  parameter HSTART  = 30  ;
  parameter VSTART  = 30  ;
  parameter HSIZE   = 1920;
  parameter VSIZE   = 1080;
  parameter CLK_DIV = 3;
`elsif TEST_PAT0
  parameter HTOTAL  = 28;
  parameter VTOTAL  = 28;
  parameter HSTART  = 10;
  parameter VSTART  = 10;
  parameter HSIZE   = 8 ;
  parameter VSIZE   = 8 ;
  parameter CLK_DIV = 1 ;
`elsif TEST_PAT1
  parameter HTOTAL  = 120;
  parameter VTOTAL  = 100;
  parameter HSTART  = 10;
  parameter VSTART  = 10;
  parameter HSIZE   = 99;
  parameter VSIZE   = 80;
  parameter CLK_DIV = 1 ;
`elsif TEST_PAT2
  parameter HTOTAL  = 1300;
  parameter VTOTAL  = 800;
  parameter HSTART  = 10;
  parameter VSTART  = 10;
  parameter HSIZE   = 1280;
  parameter VSIZE   = 720;
  parameter CLK_DIV = 1 ;
`elsif TEST_PAT3
  parameter HTOTAL  = 850;
  parameter VTOTAL  = 650;
  parameter HSTART  = 10;
  parameter VSTART  = 10;
  parameter HSIZE   = 800;
  parameter VSIZE   = 600;
  parameter CLK_DIV = 1 ;
`endif

  always @(posedge clk or negedge rstn) begin
      if (~rstn) begin
          clk_div <= `DLY 0;
      end
      else if (clk_div == (CLK_DIV - 1)) begin
          clk_div <= `DLY 0;
      end
      else begin
          clk_div <= `DLY clk_div + 1;
      end
  end

  always @(posedge clk or negedge rstn) begin
      if (~rstn) begin
          hcnt <= `DLY 0;
      end
      else if (clk_div == (CLK_DIV - 1)) begin
          if (hcnt == (HTOTAL - 1)) begin
              hcnt <= `DLY 0;
          end
          else begin
              hcnt <= `DLY hcnt + 1;
          end
      end
  end

  always @(posedge clk or negedge rstn) begin
      if (~rstn) begin
          vcnt <= `DLY 0;
      end
      else if (clk_div == (CLK_DIV - 1)) begin
          if ((hcnt == (HTOTAL - 1)) & (vcnt == (VTOTAL - 1))) begin
              vcnt <= `DLY 0;
          end
          else if (hcnt == (HTOTAL - 1))begin
              vcnt <= `DLY vcnt + 1;
          end
      end
  end

  assign pic_dat_en = (hcnt >= (HSTART        )) &
                      (hcnt <  (HSTART + HSIZE)) &
                      (vcnt >= (VSTART        )) &
                      (vcnt <  (VSTART + VSIZE)) &
                      (clk_div == (CLK_DIV - 1)) ;

  assign pic_addr = (vcnt - VSTART) * HSIZE + (hcnt - HSTART);

`ifdef SIMULATION
  initial begin
      $readmemh("bmp_data.txt", bmp_data_mem);
  end

  assign pic_data = pic_dat_en ? bmp_data_mem[(vcnt - VSTART) * HSIZE + (hcnt - HSTART)] : 24'h0;
`elsif TEST_PAT0
  always @(*) begin
      case (pic_addr)
          6'h00  : pic_data = 24'h0900b2;
          6'h01  : pic_data = 24'h330099;
          6'h02  : pic_data = 24'h600073;
          6'h03  : pic_data = 24'h8b0054;
          6'h04  : pic_data = 24'hb70034;
          6'h05  : pic_data = 24'he20015;
          6'h06  : pic_data = 24'hff0f00;
          6'h07  : pic_data = 24'hff3b00;
          6'h08  : pic_data = 24'h330099;
          6'h09  : pic_data = 24'h600073;
          6'h0A  : pic_data = 24'h8b0054;
          6'h0B  : pic_data = 24'hb70034;
          6'h0C  : pic_data = 24'he20015;
          6'h0D  : pic_data = 24'hff0f00;
          6'h0E  : pic_data = 24'hff3b00;
          6'h0F  : pic_data = 24'hff6600;
          6'h10  : pic_data = 24'h600073;
          6'h11  : pic_data = 24'h8b0054;
          6'h12  : pic_data = 24'hb70034;
          6'h13  : pic_data = 24'he20015;
          6'h14  : pic_data = 24'hff0f00;
          6'h15  : pic_data = 24'hff3b00;
          6'h16  : pic_data = 24'hff6600;
          6'h17  : pic_data = 24'hff9900;
          6'h18  : pic_data = 24'h8b0054;
          6'h19  : pic_data = 24'hb70034;
          6'h1A  : pic_data = 24'he20015;
          6'h1B  : pic_data = 24'hff0f00;
          6'h1C  : pic_data = 24'hff3b00;
          6'h1D  : pic_data = 24'hff6600;
          6'h1E  : pic_data = 24'hff9900;
          6'h1F  : pic_data = 24'hffc100;
          6'h20  : pic_data = 24'hb70034;
          6'h21  : pic_data = 24'he20015;
          6'h22  : pic_data = 24'hff0f00;
          6'h23  : pic_data = 24'hff3b00;
          6'h24  : pic_data = 24'hff6600;
          6'h25  : pic_data = 24'hff9900;
          6'h26  : pic_data = 24'hffc100;
          6'h27  : pic_data = 24'hffed00;
          6'h28  : pic_data = 24'he20015;
          6'h29  : pic_data = 24'hff0f00;
          6'h2A  : pic_data = 24'hff3b00;
          6'h2B  : pic_data = 24'hff6600;
          6'h2C  : pic_data = 24'hff9900;
          6'h2D  : pic_data = 24'hffc100;
          6'h2E  : pic_data = 24'hffed00;
          6'h2F  : pic_data = 24'hffff00;
          6'h30  : pic_data = 24'hff0f00;
          6'h31  : pic_data = 24'hff3b00;
          6'h32  : pic_data = 24'hff6600;
          6'h33  : pic_data = 24'hff9900;
          6'h34  : pic_data = 24'hffc100;
          6'h35  : pic_data = 24'hffed00;
          6'h36  : pic_data = 24'hffff00;
          6'h37  : pic_data = 24'hffff00;
          6'h38  : pic_data = 24'hff3b00;
          6'h39  : pic_data = 24'hff6600;
          6'h3A  : pic_data = 24'hff9900;
          6'h3B  : pic_data = 24'hffc100;
          6'h3C  : pic_data = 24'hffed00;
          6'h3D  : pic_data = 24'hffff00;
          6'h3E  : pic_data = 24'hffff00;
          default: pic_data = 24'hffff00;
      endcase
  end
`elsif TEST_PAT1
  always @(*) begin
      case (pic_addr)
          13'h0000 : pic_data = 24'hff0000;
          13'h0001 : pic_data = 24'hff0d00;
          13'h0002 : pic_data = 24'hff1800;
          13'h0003 : pic_data = 24'hff3400;
          13'h0004 : pic_data = 24'hff3e00;
          13'h0005 : pic_data = 24'hff4d00;
          13'h0006 : pic_data = 24'hff5800;
          13'h0007 : pic_data = 24'hff6400;
          13'h0008 : pic_data = 24'hff8000;
          13'h0009 : pic_data = 24'hff8a00;
          13'h000A : pic_data = 24'hff9900;
          13'h000B : pic_data = 24'hffa300;
          13'h000C : pic_data = 24'hffb200;
          13'h000D : pic_data = 24'hffcb00;
          13'h000E : pic_data = 24'hffd600;
          13'h000F : pic_data = 24'hffe600;
          13'h0010 : pic_data = 24'hffef00;
          13'h0011 : pic_data = 24'hffff00;
          13'h0012 : pic_data = 24'he6ff00;
          13'h0013 : pic_data = 24'hdcff00;
          13'h0014 : pic_data = 24'hccff00;
          13'h0015 : pic_data = 24'hb3ff00;
          13'h0016 : pic_data = 24'hb5ff00;
          13'h0017 : pic_data = 24'h9aff00;
          13'h0018 : pic_data = 24'h90ff00;
          13'h0019 : pic_data = 24'h80ff00;
          13'h001A : pic_data = 24'h66ff00;
          13'h001B : pic_data = 24'h68ff00;
          13'h001C : pic_data = 24'h50ff00;
          13'h001D : pic_data = 24'h44ff00;
          13'h001E : pic_data = 24'h33ff00;
          13'h001F : pic_data = 24'h1bff00;
          13'h0020 : pic_data = 24'h1cff00;
          13'h0021 : pic_data = 24'h01ff00;
          13'h0022 : pic_data = 24'h00ff06;
          13'h0023 : pic_data = 24'h00ff19;
          13'h0024 : pic_data = 24'h00ff2e;
          13'h0025 : pic_data = 24'h00ff3a;
          13'h0026 : pic_data = 24'h00ff4e;
          13'h0027 : pic_data = 24'h00ff52;
          13'h0028 : pic_data = 24'h00ff65;
          13'h0029 : pic_data = 24'h00ff7c;
          13'h002A : pic_data = 24'h00ff86;
          13'h002B : pic_data = 24'h00ff9a;
          13'h002C : pic_data = 24'h00ff9e;
          13'h002D : pic_data = 24'h00ffb3;
          13'h002E : pic_data = 24'h00ffc6;
          13'h002F : pic_data = 24'h00ffd2;
          13'h0030 : pic_data = 24'h00ffe7;
          13'h0031 : pic_data = 24'h00ffea;
          13'h0032 : pic_data = 24'h00ffff;
          13'h0033 : pic_data = 24'h00ebff;
          13'h0034 : pic_data = 24'h00e1ff;
          13'h0035 : pic_data = 24'h00cbff;
          13'h0036 : pic_data = 24'h00b8ff;
          13'h0037 : pic_data = 24'h00b4ff;
          13'h0038 : pic_data = 24'h009fff;
          13'h0039 : pic_data = 24'h0095ff;
          13'h003A : pic_data = 24'h007fff;
          13'h003B : pic_data = 24'h006cff;
          13'h003C : pic_data = 24'h0067ff;
          13'h003D : pic_data = 24'h0054ff;
          13'h003E : pic_data = 24'h0049ff;
          13'h003F : pic_data = 24'h0032ff;
          13'h0040 : pic_data = 24'h0020ff;
          13'h0041 : pic_data = 24'h001bff;
          13'h0042 : pic_data = 24'h0008ff;
          13'h0043 : pic_data = 24'h0100ff;
          13'h0044 : pic_data = 24'h1a00ff;
          13'h0045 : pic_data = 24'h2a00ff;
          13'h0046 : pic_data = 24'h3500ff;
          13'h0047 : pic_data = 24'h4f00ff;
          13'h0048 : pic_data = 24'h4d00ff;
          13'h0049 : pic_data = 24'h6600ff;
          13'h004A : pic_data = 24'h7600ff;
          13'h004B : pic_data = 24'h8100ff;
          13'h004C : pic_data = 24'h9b00ff;
          13'h004D : pic_data = 24'h9900ff;
          13'h004E : pic_data = 24'hb400ff;
          13'h004F : pic_data = 24'hc200ff;
          13'h0050 : pic_data = 24'hcc00ff;
          13'h0051 : pic_data = 24'he800ff;
          13'h0052 : pic_data = 24'he500ff;
          13'h0053 : pic_data = 24'hff00ff;
          13'h0054 : pic_data = 24'hff00f0;
          13'h0055 : pic_data = 24'hff00e5;
          13'h0056 : pic_data = 24'hff00ca;
          13'h0057 : pic_data = 24'hff00bd;
          13'h0058 : pic_data = 24'hff00b3;
          13'h0059 : pic_data = 24'hff00a4;
          13'h005A : pic_data = 24'hff0099;
          13'h005B : pic_data = 24'hff007e;
          13'h005C : pic_data = 24'hff0071;
          13'h005D : pic_data = 24'hff0066;
          13'h005E : pic_data = 24'hff0058;
          13'h005F : pic_data = 24'hff004e;
          13'h0060 : pic_data = 24'hff0031;
          13'h0061 : pic_data = 24'hff0025;
          13'h0062 : pic_data = 24'hff0018;
          13'h0063 : pic_data = 24'hff0000;
          13'h0064 : pic_data = 24'hff0c00;
          13'h0065 : pic_data = 24'hff1800;
          13'h0066 : pic_data = 24'hff3400;
          13'h0067 : pic_data = 24'hff3e00;
          13'h0068 : pic_data = 24'hff4d00;
          13'h0069 : pic_data = 24'hff5800;
          13'h006A : pic_data = 24'hff6400;
          13'h006B : pic_data = 24'hff8000;
          13'h006C : pic_data = 24'hff8a00;
          13'h006D : pic_data = 24'hff9900;
          13'h006E : pic_data = 24'hffa300;
          13'h006F : pic_data = 24'hffb200;
          13'h0070 : pic_data = 24'hffcb00;
          13'h0071 : pic_data = 24'hffd600;
          13'h0072 : pic_data = 24'hffe600;
          13'h0073 : pic_data = 24'hffef00;
          13'h0074 : pic_data = 24'hffff00;
          13'h0075 : pic_data = 24'he6ff00;
          13'h0076 : pic_data = 24'hdcff00;
          13'h0077 : pic_data = 24'hccff00;
          13'h0078 : pic_data = 24'hb3ff00;
          13'h0079 : pic_data = 24'hb5ff00;
          13'h007A : pic_data = 24'h9aff00;
          13'h007B : pic_data = 24'h90ff00;
          13'h007C : pic_data = 24'h80ff00;
          13'h007D : pic_data = 24'h66ff00;
          13'h007E : pic_data = 24'h68ff00;
          13'h007F : pic_data = 24'h4fff00;
          13'h0080 : pic_data = 24'h44ff00;
          13'h0081 : pic_data = 24'h33ff00;
          13'h0082 : pic_data = 24'h1bff00;
          13'h0083 : pic_data = 24'h1cff00;
          13'h0084 : pic_data = 24'h01ff00;
          13'h0085 : pic_data = 24'h00ff06;
          13'h0086 : pic_data = 24'h00ff19;
          13'h0087 : pic_data = 24'h00ff2e;
          13'h0088 : pic_data = 24'h00ff3a;
          13'h0089 : pic_data = 24'h00ff4e;
          13'h008A : pic_data = 24'h00ff52;
          13'h008B : pic_data = 24'h00ff65;
          13'h008C : pic_data = 24'h00ff7c;
          13'h008D : pic_data = 24'h00ff86;
          13'h008E : pic_data = 24'h00ff9a;
          13'h008F : pic_data = 24'h00ff9e;
          13'h0090 : pic_data = 24'h00ffb3;
          13'h0091 : pic_data = 24'h00ffc6;
          13'h0092 : pic_data = 24'h00ffd2;
          13'h0093 : pic_data = 24'h00ffe7;
          13'h0094 : pic_data = 24'h00ffea;
          13'h0095 : pic_data = 24'h00ffff;
          13'h0096 : pic_data = 24'h00ebff;
          13'h0097 : pic_data = 24'h00e1ff;
          13'h0098 : pic_data = 24'h00cbff;
          13'h0099 : pic_data = 24'h00b8ff;
          13'h009A : pic_data = 24'h00b4ff;
          13'h009B : pic_data = 24'h009fff;
          13'h009C : pic_data = 24'h0095ff;
          13'h009D : pic_data = 24'h007fff;
          13'h009E : pic_data = 24'h006cff;
          13'h009F : pic_data = 24'h0067ff;
          13'h00A0 : pic_data = 24'h0054ff;
          13'h00A1 : pic_data = 24'h0048ff;
          13'h00A2 : pic_data = 24'h0032ff;
          13'h00A3 : pic_data = 24'h0020ff;
          13'h00A4 : pic_data = 24'h001aff;
          13'h00A5 : pic_data = 24'h0007ff;
          13'h00A6 : pic_data = 24'h0100ff;
          13'h00A7 : pic_data = 24'h1a00ff;
          13'h00A8 : pic_data = 24'h2a00ff;
          13'h00A9 : pic_data = 24'h3500ff;
          13'h00AA : pic_data = 24'h4f00ff;
          13'h00AB : pic_data = 24'h4d00ff;
          13'h00AC : pic_data = 24'h6600ff;
          13'h00AD : pic_data = 24'h7600ff;
          13'h00AE : pic_data = 24'h8100ff;
          13'h00AF : pic_data = 24'h9b00ff;
          13'h00B0 : pic_data = 24'h9900ff;
          13'h00B1 : pic_data = 24'hb400ff;
          13'h00B2 : pic_data = 24'hc200ff;
          13'h00B3 : pic_data = 24'hcc00ff;
          13'h00B4 : pic_data = 24'he800ff;
          13'h00B5 : pic_data = 24'he500ff;
          13'h00B6 : pic_data = 24'hff00ff;
          13'h00B7 : pic_data = 24'hff00f1;
          13'h00B8 : pic_data = 24'hff00e5;
          13'h00B9 : pic_data = 24'hff00ca;
          13'h00BA : pic_data = 24'hff00bd;
          13'h00BB : pic_data = 24'hff00b3;
          13'h00BC : pic_data = 24'hff00a4;
          13'h00BD : pic_data = 24'hff0099;
          13'h00BE : pic_data = 24'hff007e;
          13'h00BF : pic_data = 24'hff0071;
          13'h00C0 : pic_data = 24'hff0066;
          13'h00C1 : pic_data = 24'hff0058;
          13'h00C2 : pic_data = 24'hff004e;
          13'h00C3 : pic_data = 24'hff0031;
          13'h00C4 : pic_data = 24'hff0025;
          13'h00C5 : pic_data = 24'hff0018;
          13'h00C6 : pic_data = 24'hfd0001;
          13'h00C7 : pic_data = 24'hfd0e01;
          13'h00C8 : pic_data = 24'hfd1a01;
          13'h00C9 : pic_data = 24'hfd3501;
          13'h00CA : pic_data = 24'hfd3f01;
          13'h00CB : pic_data = 24'hfd4e01;
          13'h00CC : pic_data = 24'hfd5901;
          13'h00CD : pic_data = 24'hfd6501;
          13'h00CE : pic_data = 24'hfd8001;
          13'h00CF : pic_data = 24'hfd8a01;
          13'h00D0 : pic_data = 24'hfd9801;
          13'h00D1 : pic_data = 24'hfda301;
          13'h00D2 : pic_data = 24'hfdb001;
          13'h00D3 : pic_data = 24'hfdca01;
          13'h00D4 : pic_data = 24'hfdd501;
          13'h00D5 : pic_data = 24'hfde401;
          13'h00D6 : pic_data = 24'hfded01;
          13'h00D7 : pic_data = 24'hfffe01;
          13'h00D8 : pic_data = 24'he4fd01;
          13'h00D9 : pic_data = 24'hdafd01;
          13'h00DA : pic_data = 24'hcbfd01;
          13'h00DB : pic_data = 24'hb2fd01;
          13'h00DC : pic_data = 24'hb3fd01;
          13'h00DD : pic_data = 24'h9afd01;
          13'h00DE : pic_data = 24'h8ffd01;
          13'h00DF : pic_data = 24'h80fd01;
          13'h00E0 : pic_data = 24'h67fd01;
          13'h00E1 : pic_data = 24'h68fd01;
          13'h00E2 : pic_data = 24'h50fd01;
          13'h00E3 : pic_data = 24'h45fd01;
          13'h00E4 : pic_data = 24'h34fd01;
          13'h00E5 : pic_data = 24'h1dfd01;
          13'h00E6 : pic_data = 24'h1dfd01;
          13'h00E7 : pic_data = 24'h03fd00;
          13'h00E8 : pic_data = 24'h01fd08;
          13'h00E9 : pic_data = 24'h01fd1b;
          13'h00EA : pic_data = 24'h01fd30;
          13'h00EB : pic_data = 24'h01fd3b;
          13'h00EC : pic_data = 24'h01fd4f;
          13'h00ED : pic_data = 24'h01fd53;
          13'h00EE : pic_data = 24'h01fd66;
          13'h00EF : pic_data = 24'h01fd7c;
          13'h00F0 : pic_data = 24'h01fd86;
          13'h00F1 : pic_data = 24'h01fd99;
          13'h00F2 : pic_data = 24'h01fd9e;
          13'h00F3 : pic_data = 24'h01fdb1;
          13'h00F4 : pic_data = 24'h01fdc5;
          13'h00F5 : pic_data = 24'h01fdd0;
          13'h00F6 : pic_data = 24'h01fde5;
          13'h00F7 : pic_data = 24'h01fde8;
          13'h00F8 : pic_data = 24'h01ffff;
          13'h00F9 : pic_data = 24'h01e9fd;
          13'h00FA : pic_data = 24'h01defd;
          13'h00FB : pic_data = 24'h01cafd;
          13'h00FC : pic_data = 24'h01b7fd;
          13'h00FD : pic_data = 24'h01b2fd;
          13'h00FE : pic_data = 24'h019efd;
          13'h00FF : pic_data = 24'h0194fd;
          13'h0100 : pic_data = 24'h017ffd;
          13'h0101 : pic_data = 24'h016cfd;
          13'h0102 : pic_data = 24'h0167fd;
          13'h0103 : pic_data = 24'h0154fd;
          13'h0104 : pic_data = 24'h014afd;
          13'h0105 : pic_data = 24'h0133fd;
          13'h0106 : pic_data = 24'h0122fd;
          13'h0107 : pic_data = 24'h011cfd;
          13'h0108 : pic_data = 24'h0109fd;
          13'h0109 : pic_data = 24'h0300fd;
          13'h010A : pic_data = 24'h1c01fd;
          13'h010B : pic_data = 24'h2b01fd;
          13'h010C : pic_data = 24'h3601fd;
          13'h010D : pic_data = 24'h5001fd;
          13'h010E : pic_data = 24'h4e01fd;
          13'h010F : pic_data = 24'h6701fd;
          13'h0110 : pic_data = 24'h7601fd;
          13'h0111 : pic_data = 24'h8101fd;
          13'h0112 : pic_data = 24'h9a01fd;
          13'h0113 : pic_data = 24'h9901fd;
          13'h0114 : pic_data = 24'hb201fd;
          13'h0115 : pic_data = 24'hc101fd;
          13'h0116 : pic_data = 24'hcb01fd;
          13'h0117 : pic_data = 24'he601fd;
          13'h0118 : pic_data = 24'he301fd;
          13'h0119 : pic_data = 24'hff01fe;
          13'h011A : pic_data = 24'hfd01ee;
          13'h011B : pic_data = 24'hfd01e3;
          13'h011C : pic_data = 24'hfd01c9;
          13'h011D : pic_data = 24'hfd01bc;
          13'h011E : pic_data = 24'hfd01b1;
          13'h011F : pic_data = 24'hfd01a3;
          13'h0120 : pic_data = 24'hfd0198;
          13'h0121 : pic_data = 24'hfd017e;
          13'h0122 : pic_data = 24'hfd0172;
          13'h0123 : pic_data = 24'hfd0166;
          13'h0124 : pic_data = 24'hfd0159;
          13'h0125 : pic_data = 24'hfd014f;
          13'h0126 : pic_data = 24'hfd0132;
          13'h0127 : pic_data = 24'hfd0127;
          13'h0128 : pic_data = 24'hfd0119;
          13'h0129 : pic_data = 24'hfa0204;
          13'h012A : pic_data = 24'hfa1004;
          13'h012B : pic_data = 24'hfa1b04;
          13'h012C : pic_data = 24'hfa3604;
          13'h012D : pic_data = 24'hfa4004;
          13'h012E : pic_data = 24'hfa4f04;
          13'h012F : pic_data = 24'hfa5904;
          13'h0130 : pic_data = 24'hfa6504;
          13'h0131 : pic_data = 24'hfa8004;
          13'h0132 : pic_data = 24'hfa8a04;
          13'h0133 : pic_data = 24'hfa9804;
          13'h0134 : pic_data = 24'hfaa204;
          13'h0135 : pic_data = 24'hfaae04;
          13'h0136 : pic_data = 24'hfac904;
          13'h0137 : pic_data = 24'hfad304;
          13'h0138 : pic_data = 24'hfae204;
          13'h0139 : pic_data = 24'hfaeb04;
          13'h013A : pic_data = 24'hfdfc04;
          13'h013B : pic_data = 24'he2fa04;
          13'h013C : pic_data = 24'hd7fa04;
          13'h013D : pic_data = 24'hcafa04;
          13'h013E : pic_data = 24'hb0fa04;
          13'h013F : pic_data = 24'hb2fa04;
          13'h0140 : pic_data = 24'h99fa04;
          13'h0141 : pic_data = 24'h8ffa04;
          13'h0142 : pic_data = 24'h80fa04;
          13'h0143 : pic_data = 24'h67fa04;
          13'h0144 : pic_data = 24'h69fa04;
          13'h0145 : pic_data = 24'h50fa04;
          13'h0146 : pic_data = 24'h46fa04;
          13'h0147 : pic_data = 24'h35fa04;
          13'h0148 : pic_data = 24'h1ffa04;
          13'h0149 : pic_data = 24'h1ffa04;
          13'h014A : pic_data = 24'h06fa03;
          13'h014B : pic_data = 24'h03fa0b;
          13'h014C : pic_data = 24'h04fa1c;
          13'h014D : pic_data = 24'h04fa32;
          13'h014E : pic_data = 24'h04fa3c;
          13'h014F : pic_data = 24'h04fa50;
          13'h0150 : pic_data = 24'h04fa54;
          13'h0151 : pic_data = 24'h04fa66;
          13'h0152 : pic_data = 24'h04fa7c;
          13'h0153 : pic_data = 24'h04fa86;
          13'h0154 : pic_data = 24'h04fa99;
          13'h0155 : pic_data = 24'h04fa9d;
          13'h0156 : pic_data = 24'h04faaf;
          13'h0157 : pic_data = 24'h04fac4;
          13'h0158 : pic_data = 24'h04facf;
          13'h0159 : pic_data = 24'h04fae3;
          13'h015A : pic_data = 24'h04fae6;
          13'h015B : pic_data = 24'h04fdfd;
          13'h015C : pic_data = 24'h04e6fa;
          13'h015D : pic_data = 24'h04dcfa;
          13'h015E : pic_data = 24'h04c9fa;
          13'h015F : pic_data = 24'h04b5fa;
          13'h0160 : pic_data = 24'h04b1fa;
          13'h0161 : pic_data = 24'h049efa;
          13'h0162 : pic_data = 24'h0493fa;
          13'h0163 : pic_data = 24'h047ffa;
          13'h0164 : pic_data = 24'h046cfa;
          13'h0165 : pic_data = 24'h0468fa;
          13'h0166 : pic_data = 24'h0455fa;
          13'h0167 : pic_data = 24'h044bfa;
          13'h0168 : pic_data = 24'h0434fa;
          13'h0169 : pic_data = 24'h0424fa;
          13'h016A : pic_data = 24'h041efa;
          13'h016B : pic_data = 24'h030bfa;
          13'h016C : pic_data = 24'h0603fa;
          13'h016D : pic_data = 24'h1d04fa;
          13'h016E : pic_data = 24'h2d04fa;
          13'h016F : pic_data = 24'h3704fa;
          13'h0170 : pic_data = 24'h5104fa;
          13'h0171 : pic_data = 24'h4f04fa;
          13'h0172 : pic_data = 24'h6704fa;
          13'h0173 : pic_data = 24'h7704fa;
          13'h0174 : pic_data = 24'h8104fa;
          13'h0175 : pic_data = 24'h9a04fa;
          13'h0176 : pic_data = 24'h9804fa;
          13'h0177 : pic_data = 24'hb004fa;
          13'h0178 : pic_data = 24'hc004fa;
          13'h0179 : pic_data = 24'hca04fa;
          13'h017A : pic_data = 24'he404fa;
          13'h017B : pic_data = 24'he104fa;
          13'h017C : pic_data = 24'hfd04fc;
          13'h017D : pic_data = 24'hfa04ec;
          13'h017E : pic_data = 24'hfa04e0;
          13'h017F : pic_data = 24'hfa04c8;
          13'h0180 : pic_data = 24'hfa04ba;
          13'h0181 : pic_data = 24'hfa04b0;
          13'h0182 : pic_data = 24'hfa04a2;
          13'h0183 : pic_data = 24'hfa0498;
          13'h0184 : pic_data = 24'hfa047e;
          13'h0185 : pic_data = 24'hfa0472;
          13'h0186 : pic_data = 24'hfa0467;
          13'h0187 : pic_data = 24'hfa0459;
          13'h0188 : pic_data = 24'hfa0451;
          13'h0189 : pic_data = 24'hfa0433;
          13'h018A : pic_data = 24'hfa0429;
          13'h018B : pic_data = 24'hfa041b;
          13'h018C : pic_data = 24'hfb0203;
          13'h018D : pic_data = 24'hfb0f03;
          13'h018E : pic_data = 24'hfb1b03;
          13'h018F : pic_data = 24'hfb3603;
          13'h0190 : pic_data = 24'hfb4003;
          13'h0191 : pic_data = 24'hfb4f03;
          13'h0192 : pic_data = 24'hfb5903;
          13'h0193 : pic_data = 24'hfb6503;
          13'h0194 : pic_data = 24'hfb8003;
          13'h0195 : pic_data = 24'hfb8a03;
          13'h0196 : pic_data = 24'hfb9803;
          13'h0197 : pic_data = 24'hfba203;
          13'h0198 : pic_data = 24'hfbae03;
          13'h0199 : pic_data = 24'hfbc903;
          13'h019A : pic_data = 24'hfbd303;
          13'h019B : pic_data = 24'hfbe203;
          13'h019C : pic_data = 24'hfbeb03;
          13'h019D : pic_data = 24'hfefd03;
          13'h019E : pic_data = 24'he2fb03;
          13'h019F : pic_data = 24'hd8fb03;
          13'h01A0 : pic_data = 24'hcbfb03;
          13'h01A1 : pic_data = 24'hb0fb03;
          13'h01A2 : pic_data = 24'hb2fb03;
          13'h01A3 : pic_data = 24'h99fb03;
          13'h01A4 : pic_data = 24'h8ffb03;
          13'h01A5 : pic_data = 24'h80fb03;
          13'h01A6 : pic_data = 24'h67fb03;
          13'h01A7 : pic_data = 24'h69fb03;
          13'h01A8 : pic_data = 24'h50fb03;
          13'h01A9 : pic_data = 24'h46fb03;
          13'h01AA : pic_data = 24'h35fb03;
          13'h01AB : pic_data = 24'h1efb03;
          13'h01AC : pic_data = 24'h1efb03;
          13'h01AD : pic_data = 24'h05fb02;
          13'h01AE : pic_data = 24'h03fb0a;
          13'h01AF : pic_data = 24'h03fb1c;
          13'h01B0 : pic_data = 24'h03fb31;
          13'h01B1 : pic_data = 24'h03fb3c;
          13'h01B2 : pic_data = 24'h03fb50;
          13'h01B3 : pic_data = 24'h03fb54;
          13'h01B4 : pic_data = 24'h03fb66;
          13'h01B5 : pic_data = 24'h03fb7c;
          13'h01B6 : pic_data = 24'h03fb86;
          13'h01B7 : pic_data = 24'h03fb99;
          13'h01B8 : pic_data = 24'h03fb9d;
          13'h01B9 : pic_data = 24'h03fbaf;
          13'h01BA : pic_data = 24'h03fbc5;
          13'h01BB : pic_data = 24'h03fbcf;
          13'h01BC : pic_data = 24'h03fbe3;
          13'h01BD : pic_data = 24'h03fbe6;
          13'h01BE : pic_data = 24'h03fdfd;
          13'h01BF : pic_data = 24'h03e7fb;
          13'h01C0 : pic_data = 24'h03dcfb;
          13'h01C1 : pic_data = 24'h03cafb;
          13'h01C2 : pic_data = 24'h03b5fb;
          13'h01C3 : pic_data = 24'h03b1fb;
          13'h01C4 : pic_data = 24'h039efb;
          13'h01C5 : pic_data = 24'h0393fb;
          13'h01C6 : pic_data = 24'h037ffb;
          13'h01C7 : pic_data = 24'h036cfb;
          13'h01C8 : pic_data = 24'h0368fb;
          13'h01C9 : pic_data = 24'h0355fb;
          13'h01CA : pic_data = 24'h034bfb;
          13'h01CB : pic_data = 24'h0334fb;
          13'h01CC : pic_data = 24'h0323fb;
          13'h01CD : pic_data = 24'h031dfb;
          13'h01CE : pic_data = 24'h030afb;
          13'h01CF : pic_data = 24'h0502fb;
          13'h01D0 : pic_data = 24'h1d03fb;
          13'h01D1 : pic_data = 24'h2d03fb;
          13'h01D2 : pic_data = 24'h3703fb;
          13'h01D3 : pic_data = 24'h5103fb;
          13'h01D4 : pic_data = 24'h4f03fb;
          13'h01D5 : pic_data = 24'h6703fb;
          13'h01D6 : pic_data = 24'h7703fb;
          13'h01D7 : pic_data = 24'h8103fb;
          13'h01D8 : pic_data = 24'h9a03fb;
          13'h01D9 : pic_data = 24'h9803fb;
          13'h01DA : pic_data = 24'hb003fb;
          13'h01DB : pic_data = 24'hc003fb;
          13'h01DC : pic_data = 24'hca03fb;
          13'h01DD : pic_data = 24'he403fb;
          13'h01DE : pic_data = 24'he103fb;
          13'h01DF : pic_data = 24'hfe03fc;
          13'h01E0 : pic_data = 24'hfb03ed;
          13'h01E1 : pic_data = 24'hfb03e1;
          13'h01E2 : pic_data = 24'hfb03c9;
          13'h01E3 : pic_data = 24'hfb03ba;
          13'h01E4 : pic_data = 24'hfb03b0;
          13'h01E5 : pic_data = 24'hfb03a2;
          13'h01E6 : pic_data = 24'hfb0398;
          13'h01E7 : pic_data = 24'hfb037e;
          13'h01E8 : pic_data = 24'hfb0372;
          13'h01E9 : pic_data = 24'hfb0367;
          13'h01EA : pic_data = 24'hfb0359;
          13'h01EB : pic_data = 24'hfb0350;
          13'h01EC : pic_data = 24'hfb0333;
          13'h01ED : pic_data = 24'hfb0328;
          13'h01EE : pic_data = 24'hfb031b;
          13'h01EF : pic_data = 24'hf90406;
          13'h01F0 : pic_data = 24'hf91106;
          13'h01F1 : pic_data = 24'hf91c06;
          13'h01F2 : pic_data = 24'hf93706;
          13'h01F3 : pic_data = 24'hf94106;
          13'h01F4 : pic_data = 24'hf94f06;
          13'h01F5 : pic_data = 24'hf95a06;
          13'h01F6 : pic_data = 24'hf96606;
          13'h01F7 : pic_data = 24'hf98006;
          13'h01F8 : pic_data = 24'hf98a06;
          13'h01F9 : pic_data = 24'hf99706;
          13'h01FA : pic_data = 24'hf9a206;
          13'h01FB : pic_data = 24'hf9ae06;
          13'h01FC : pic_data = 24'hf9c806;
          13'h01FD : pic_data = 24'hf9d206;
          13'h01FE : pic_data = 24'hf9e106;
          13'h01FF : pic_data = 24'hf9ea06;
          13'h0200 : pic_data = 24'hfbfa06;
          13'h0201 : pic_data = 24'he1f906;
          13'h0202 : pic_data = 24'hd6f906;
          13'h0203 : pic_data = 24'hc9f906;
          13'h0204 : pic_data = 24'hb0f906;
          13'h0205 : pic_data = 24'hb1f906;
          13'h0206 : pic_data = 24'h99f906;
          13'h0207 : pic_data = 24'h8ef906;
          13'h0208 : pic_data = 24'h80f906;
          13'h0209 : pic_data = 24'h68f906;
          13'h020A : pic_data = 24'h69f906;
          13'h020B : pic_data = 24'h51f906;
          13'h020C : pic_data = 24'h47f906;
          13'h020D : pic_data = 24'h36f906;
          13'h020E : pic_data = 24'h20f906;
          13'h020F : pic_data = 24'h20f906;
          13'h0210 : pic_data = 24'h08f905;
          13'h0211 : pic_data = 24'h05f90c;
          13'h0212 : pic_data = 24'h06f91d;
          13'h0213 : pic_data = 24'h06f933;
          13'h0214 : pic_data = 24'h06f93d;
          13'h0215 : pic_data = 24'h06f950;
          13'h0216 : pic_data = 24'h06f955;
          13'h0217 : pic_data = 24'h06f967;
          13'h0218 : pic_data = 24'h06f97b;
          13'h0219 : pic_data = 24'h06f986;
          13'h021A : pic_data = 24'h06f998;
          13'h021B : pic_data = 24'h06f99d;
          13'h021C : pic_data = 24'h06f9af;
          13'h021D : pic_data = 24'h06f9c3;
          13'h021E : pic_data = 24'h06f9cd;
          13'h021F : pic_data = 24'h06f9e2;
          13'h0220 : pic_data = 24'h06f9e5;
          13'h0221 : pic_data = 24'h06fbfb;
          13'h0222 : pic_data = 24'h06e5f9;
          13'h0223 : pic_data = 24'h06dbf9;
          13'h0224 : pic_data = 24'h06c8f9;
          13'h0225 : pic_data = 24'h06b5f9;
          13'h0226 : pic_data = 24'h06b0f9;
          13'h0227 : pic_data = 24'h069df9;
          13'h0228 : pic_data = 24'h0693f9;
          13'h0229 : pic_data = 24'h067ff9;
          13'h022A : pic_data = 24'h066df9;
          13'h022B : pic_data = 24'h0668f9;
          13'h022C : pic_data = 24'h0655f9;
          13'h022D : pic_data = 24'h064cf9;
          13'h022E : pic_data = 24'h0635f9;
          13'h022F : pic_data = 24'h0625f9;
          13'h0230 : pic_data = 24'h061ff9;
          13'h0231 : pic_data = 24'h050df9;
          13'h0232 : pic_data = 24'h0805f9;
          13'h0233 : pic_data = 24'h1e06f9;
          13'h0234 : pic_data = 24'h2e06f9;
          13'h0235 : pic_data = 24'h3806f9;
          13'h0236 : pic_data = 24'h5106f9;
          13'h0237 : pic_data = 24'h5006f9;
          13'h0238 : pic_data = 24'h6806f9;
          13'h0239 : pic_data = 24'h7706f9;
          13'h023A : pic_data = 24'h8106f9;
          13'h023B : pic_data = 24'h9906f9;
          13'h023C : pic_data = 24'h9806f9;
          13'h023D : pic_data = 24'hb006f9;
          13'h023E : pic_data = 24'hbf06f9;
          13'h023F : pic_data = 24'hc906f9;
          13'h0240 : pic_data = 24'he306f9;
          13'h0241 : pic_data = 24'he006f9;
          13'h0242 : pic_data = 24'hfb06fa;
          13'h0243 : pic_data = 24'hf906ea;
          13'h0244 : pic_data = 24'hf906df;
          13'h0245 : pic_data = 24'hf906c7;
          13'h0246 : pic_data = 24'hf906ba;
          13'h0247 : pic_data = 24'hf906af;
          13'h0248 : pic_data = 24'hf906a2;
          13'h0249 : pic_data = 24'hf90697;
          13'h024A : pic_data = 24'hf9067e;
          13'h024B : pic_data = 24'hf90672;
          13'h024C : pic_data = 24'hf90667;
          13'h024D : pic_data = 24'hf9065a;
          13'h024E : pic_data = 24'hf90651;
          13'h024F : pic_data = 24'hf90634;
          13'h0250 : pic_data = 24'hf9062a;
          13'h0251 : pic_data = 24'hf9061c;
          13'h0252 : pic_data = 24'hf60709;
          13'h0253 : pic_data = 24'hf61409;
          13'h0254 : pic_data = 24'hf61e09;
          13'h0255 : pic_data = 24'hf63909;
          13'h0256 : pic_data = 24'hf64209;
          13'h0257 : pic_data = 24'hf65009;
          13'h0258 : pic_data = 24'hf65a09;
          13'h0259 : pic_data = 24'hf66609;
          13'h025A : pic_data = 24'hf68009;
          13'h025B : pic_data = 24'hf68909;
          13'h025C : pic_data = 24'hf69709;
          13'h025D : pic_data = 24'hf6a109;
          13'h025E : pic_data = 24'hf6ad09;
          13'h025F : pic_data = 24'hf6c609;
          13'h0260 : pic_data = 24'hf6d009;
          13'h0261 : pic_data = 24'hf6df09;
          13'h0262 : pic_data = 24'hf6e809;
          13'h0263 : pic_data = 24'hf9f809;
          13'h0264 : pic_data = 24'hdff609;
          13'h0265 : pic_data = 24'hd5f609;
          13'h0266 : pic_data = 24'hc7f609;
          13'h0267 : pic_data = 24'haff609;
          13'h0268 : pic_data = 24'hb1f609;
          13'h0269 : pic_data = 24'h98f609;
          13'h026A : pic_data = 24'h8ef609;
          13'h026B : pic_data = 24'h80f609;
          13'h026C : pic_data = 24'h68f609;
          13'h026D : pic_data = 24'h6af609;
          13'h026E : pic_data = 24'h51f609;
          13'h026F : pic_data = 24'h48f609;
          13'h0270 : pic_data = 24'h38f609;
          13'h0271 : pic_data = 24'h22f609;
          13'h0272 : pic_data = 24'h22f609;
          13'h0273 : pic_data = 24'h0bf608;
          13'h0274 : pic_data = 24'h08f60f;
          13'h0275 : pic_data = 24'h09f61f;
          13'h0276 : pic_data = 24'h09f635;
          13'h0277 : pic_data = 24'h09f63e;
          13'h0278 : pic_data = 24'h09f651;
          13'h0279 : pic_data = 24'h09f655;
          13'h027A : pic_data = 24'h09f667;
          13'h027B : pic_data = 24'h09f67b;
          13'h027C : pic_data = 24'h09f686;
          13'h027D : pic_data = 24'h09f698;
          13'h027E : pic_data = 24'h09f69c;
          13'h027F : pic_data = 24'h09f6ae;
          13'h0280 : pic_data = 24'h09f6c1;
          13'h0281 : pic_data = 24'h09f6cc;
          13'h0282 : pic_data = 24'h09f6e0;
          13'h0283 : pic_data = 24'h09f6e3;
          13'h0284 : pic_data = 24'h09f8f8;
          13'h0285 : pic_data = 24'h09e4f6;
          13'h0286 : pic_data = 24'h09d9f6;
          13'h0287 : pic_data = 24'h09c6f6;
          13'h0288 : pic_data = 24'h09b4f6;
          13'h0289 : pic_data = 24'h09b0f6;
          13'h028A : pic_data = 24'h099df6;
          13'h028B : pic_data = 24'h0992f6;
          13'h028C : pic_data = 24'h097ff6;
          13'h028D : pic_data = 24'h096df6;
          13'h028E : pic_data = 24'h0969f6;
          13'h028F : pic_data = 24'h0956f6;
          13'h0290 : pic_data = 24'h094df6;
          13'h0291 : pic_data = 24'h0937f6;
          13'h0292 : pic_data = 24'h0927f6;
          13'h0293 : pic_data = 24'h0921f6;
          13'h0294 : pic_data = 24'h0810f6;
          13'h0295 : pic_data = 24'h0b08f6;
          13'h0296 : pic_data = 24'h2009f6;
          13'h0297 : pic_data = 24'h3009f6;
          13'h0298 : pic_data = 24'h3909f6;
          13'h0299 : pic_data = 24'h5209f6;
          13'h029A : pic_data = 24'h5009f6;
          13'h029B : pic_data = 24'h6809f6;
          13'h029C : pic_data = 24'h7709f6;
          13'h029D : pic_data = 24'h8209f6;
          13'h029E : pic_data = 24'h9909f6;
          13'h029F : pic_data = 24'h9709f6;
          13'h02A0 : pic_data = 24'haf09f6;
          13'h02A1 : pic_data = 24'hbd09f6;
          13'h02A2 : pic_data = 24'hc709f6;
          13'h02A3 : pic_data = 24'he109f6;
          13'h02A4 : pic_data = 24'hde09f6;
          13'h02A5 : pic_data = 24'hf909f8;
          13'h02A6 : pic_data = 24'hf609e8;
          13'h02A7 : pic_data = 24'hf609de;
          13'h02A8 : pic_data = 24'hf609c5;
          13'h02A9 : pic_data = 24'hf609b9;
          13'h02AA : pic_data = 24'hf609af;
          13'h02AB : pic_data = 24'hf609a1;
          13'h02AC : pic_data = 24'hf60997;
          13'h02AD : pic_data = 24'hf6097e;
          13'h02AE : pic_data = 24'hf60972;
          13'h02AF : pic_data = 24'hf60968;
          13'h02B0 : pic_data = 24'hf6095a;
          13'h02B1 : pic_data = 24'hf60951;
          13'h02B2 : pic_data = 24'hf60936;
          13'h02B3 : pic_data = 24'hf6092c;
          13'h02B4 : pic_data = 24'hf6091e;
          13'h02B5 : pic_data = 24'hf70708;
          13'h02B6 : pic_data = 24'hf71308;
          13'h02B7 : pic_data = 24'hf71e08;
          13'h02B8 : pic_data = 24'hf73908;
          13'h02B9 : pic_data = 24'hf74208;
          13'h02BA : pic_data = 24'hf75008;
          13'h02BB : pic_data = 24'hf75a08;
          13'h02BC : pic_data = 24'hf76608;
          13'h02BD : pic_data = 24'hf78008;
          13'h02BE : pic_data = 24'hf78908;
          13'h02BF : pic_data = 24'hf79708;
          13'h02C0 : pic_data = 24'hf7a108;
          13'h02C1 : pic_data = 24'hf7ad08;
          13'h02C2 : pic_data = 24'hf7c608;
          13'h02C3 : pic_data = 24'hf7d008;
          13'h02C4 : pic_data = 24'hf7df08;
          13'h02C5 : pic_data = 24'hf7e808;
          13'h02C6 : pic_data = 24'hfaf908;
          13'h02C7 : pic_data = 24'hdff708;
          13'h02C8 : pic_data = 24'hd5f708;
          13'h02C9 : pic_data = 24'hc7f708;
          13'h02CA : pic_data = 24'haff708;
          13'h02CB : pic_data = 24'hb1f708;
          13'h02CC : pic_data = 24'h98f708;
          13'h02CD : pic_data = 24'h8ef708;
          13'h02CE : pic_data = 24'h80f708;
          13'h02CF : pic_data = 24'h68f708;
          13'h02D0 : pic_data = 24'h6af708;
          13'h02D1 : pic_data = 24'h51f708;
          13'h02D2 : pic_data = 24'h48f708;
          13'h02D3 : pic_data = 24'h38f708;
          13'h02D4 : pic_data = 24'h21f708;
          13'h02D5 : pic_data = 24'h21f708;
          13'h02D6 : pic_data = 24'h0af707;
          13'h02D7 : pic_data = 24'h08f70e;
          13'h02D8 : pic_data = 24'h08f71f;
          13'h02D9 : pic_data = 24'h08f735;
          13'h02DA : pic_data = 24'h08f73e;
          13'h02DB : pic_data = 24'h08f751;
          13'h02DC : pic_data = 24'h08f755;
          13'h02DD : pic_data = 24'h08f767;
          13'h02DE : pic_data = 24'h08f77b;
          13'h02DF : pic_data = 24'h08f786;
          13'h02E0 : pic_data = 24'h08f798;
          13'h02E1 : pic_data = 24'h08f79c;
          13'h02E2 : pic_data = 24'h08f7ae;
          13'h02E3 : pic_data = 24'h08f7c1;
          13'h02E4 : pic_data = 24'h08f7cc;
          13'h02E5 : pic_data = 24'h08f7e0;
          13'h02E6 : pic_data = 24'h08f7e3;
          13'h02E7 : pic_data = 24'h08f9f9;
          13'h02E8 : pic_data = 24'h08e4f7;
          13'h02E9 : pic_data = 24'h08d9f7;
          13'h02EA : pic_data = 24'h08c6f7;
          13'h02EB : pic_data = 24'h08b4f7;
          13'h02EC : pic_data = 24'h08b0f7;
          13'h02ED : pic_data = 24'h089df7;
          13'h02EE : pic_data = 24'h0892f7;
          13'h02EF : pic_data = 24'h087ff7;
          13'h02F0 : pic_data = 24'h086df7;
          13'h02F1 : pic_data = 24'h0869f7;
          13'h02F2 : pic_data = 24'h0856f7;
          13'h02F3 : pic_data = 24'h084df7;
          13'h02F4 : pic_data = 24'h0837f7;
          13'h02F5 : pic_data = 24'h0826f7;
          13'h02F6 : pic_data = 24'h0820f7;
          13'h02F7 : pic_data = 24'h080ff7;
          13'h02F8 : pic_data = 24'h0a07f7;
          13'h02F9 : pic_data = 24'h2008f7;
          13'h02FA : pic_data = 24'h3008f7;
          13'h02FB : pic_data = 24'h3908f7;
          13'h02FC : pic_data = 24'h5208f7;
          13'h02FD : pic_data = 24'h5008f7;
          13'h02FE : pic_data = 24'h6808f7;
          13'h02FF : pic_data = 24'h7708f7;
          13'h0300 : pic_data = 24'h8208f7;
          13'h0301 : pic_data = 24'h9908f7;
          13'h0302 : pic_data = 24'h9708f7;
          13'h0303 : pic_data = 24'haf08f7;
          13'h0304 : pic_data = 24'hbd08f7;
          13'h0305 : pic_data = 24'hc708f7;
          13'h0306 : pic_data = 24'he108f7;
          13'h0307 : pic_data = 24'hde08f7;
          13'h0308 : pic_data = 24'hfa08f9;
          13'h0309 : pic_data = 24'hf708e8;
          13'h030A : pic_data = 24'hf708de;
          13'h030B : pic_data = 24'hf708c5;
          13'h030C : pic_data = 24'hf708b9;
          13'h030D : pic_data = 24'hf708af;
          13'h030E : pic_data = 24'hf708a1;
          13'h030F : pic_data = 24'hf70897;
          13'h0310 : pic_data = 24'hf7087e;
          13'h0311 : pic_data = 24'hf70872;
          13'h0312 : pic_data = 24'hf70868;
          13'h0313 : pic_data = 24'hf7085a;
          13'h0314 : pic_data = 24'hf70851;
          13'h0315 : pic_data = 24'hf70836;
          13'h0316 : pic_data = 24'hf7082b;
          13'h0317 : pic_data = 24'hf7081e;
          13'h0318 : pic_data = 24'hf4090a;
          13'h0319 : pic_data = 24'hf4150a;
          13'h031A : pic_data = 24'hf4200a;
          13'h031B : pic_data = 24'hf43a0a;
          13'h031C : pic_data = 24'hf4430a;
          13'h031D : pic_data = 24'hf4510a;
          13'h031E : pic_data = 24'hf45b0a;
          13'h031F : pic_data = 24'hf4660a;
          13'h0320 : pic_data = 24'hf4800a;
          13'h0321 : pic_data = 24'hf4890a;
          13'h0322 : pic_data = 24'hf4970a;
          13'h0323 : pic_data = 24'hf4a10a;
          13'h0324 : pic_data = 24'hf4ac0a;
          13'h0325 : pic_data = 24'hf4c50a;
          13'h0326 : pic_data = 24'hf4cf0a;
          13'h0327 : pic_data = 24'hf4dd0a;
          13'h0328 : pic_data = 24'hf4e60a;
          13'h0329 : pic_data = 24'hf7f60a;
          13'h032A : pic_data = 24'hdef40a;
          13'h032B : pic_data = 24'hd3f40a;
          13'h032C : pic_data = 24'hc7f40a;
          13'h032D : pic_data = 24'haef40a;
          13'h032E : pic_data = 24'hb0f40a;
          13'h032F : pic_data = 24'h98f40a;
          13'h0330 : pic_data = 24'h8ef40a;
          13'h0331 : pic_data = 24'h80f40a;
          13'h0332 : pic_data = 24'h68f40a;
          13'h0333 : pic_data = 24'h6af40a;
          13'h0334 : pic_data = 24'h52f40a;
          13'h0335 : pic_data = 24'h49f40a;
          13'h0336 : pic_data = 24'h39f40a;
          13'h0337 : pic_data = 24'h23f40a;
          13'h0338 : pic_data = 24'h23f40a;
          13'h0339 : pic_data = 24'h0cf409;
          13'h033A : pic_data = 24'h0af410;
          13'h033B : pic_data = 24'h0af421;
          13'h033C : pic_data = 24'h0af435;
          13'h033D : pic_data = 24'h0af43f;
          13'h033E : pic_data = 24'h0af452;
          13'h033F : pic_data = 24'h0af456;
          13'h0340 : pic_data = 24'h0af467;
          13'h0341 : pic_data = 24'h0af47b;
          13'h0342 : pic_data = 24'h0af486;
          13'h0343 : pic_data = 24'h0af498;
          13'h0344 : pic_data = 24'h0af49c;
          13'h0345 : pic_data = 24'h0af4ad;
          13'h0346 : pic_data = 24'h0af4c0;
          13'h0347 : pic_data = 24'h0af4cb;
          13'h0348 : pic_data = 24'h0af4de;
          13'h0349 : pic_data = 24'h0af4e1;
          13'h034A : pic_data = 24'h0af7f7;
          13'h034B : pic_data = 24'h0ae2f4;
          13'h034C : pic_data = 24'h0ad8f4;
          13'h034D : pic_data = 24'h0ac6f4;
          13'h034E : pic_data = 24'h0ab3f4;
          13'h034F : pic_data = 24'h0aaff4;
          13'h0350 : pic_data = 24'h0a9cf4;
          13'h0351 : pic_data = 24'h0a92f4;
          13'h0352 : pic_data = 24'h0a7ff4;
          13'h0353 : pic_data = 24'h0a6df4;
          13'h0354 : pic_data = 24'h0a69f4;
          13'h0355 : pic_data = 24'h0a57f4;
          13'h0356 : pic_data = 24'h0a4df4;
          13'h0357 : pic_data = 24'h0a38f4;
          13'h0358 : pic_data = 24'h0a28f4;
          13'h0359 : pic_data = 24'h0a22f4;
          13'h035A : pic_data = 24'h0a11f4;
          13'h035B : pic_data = 24'h0c09f4;
          13'h035C : pic_data = 24'h220af4;
          13'h035D : pic_data = 24'h310af4;
          13'h035E : pic_data = 24'h3a0af4;
          13'h035F : pic_data = 24'h530af4;
          13'h0360 : pic_data = 24'h510af4;
          13'h0361 : pic_data = 24'h680af4;
          13'h0362 : pic_data = 24'h770af4;
          13'h0363 : pic_data = 24'h820af4;
          13'h0364 : pic_data = 24'h990af4;
          13'h0365 : pic_data = 24'h970af4;
          13'h0366 : pic_data = 24'hae0af4;
          13'h0367 : pic_data = 24'hbc0af4;
          13'h0368 : pic_data = 24'hc60af4;
          13'h0369 : pic_data = 24'hdf0af4;
          13'h036A : pic_data = 24'hdc0af4;
          13'h036B : pic_data = 24'hf70af6;
          13'h036C : pic_data = 24'hf40ae7;
          13'h036D : pic_data = 24'hf40adc;
          13'h036E : pic_data = 24'hf40ac5;
          13'h036F : pic_data = 24'hf40ab8;
          13'h0370 : pic_data = 24'hf40aae;
          13'h0371 : pic_data = 24'hf40aa1;
          13'h0372 : pic_data = 24'hf40a97;
          13'h0373 : pic_data = 24'hf40a7e;
          13'h0374 : pic_data = 24'hf40a72;
          13'h0375 : pic_data = 24'hf40a68;
          13'h0376 : pic_data = 24'hf40a5b;
          13'h0377 : pic_data = 24'hf40a52;
          13'h0378 : pic_data = 24'hf40a37;
          13'h0379 : pic_data = 24'hf40a2d;
          13'h037A : pic_data = 24'hf40a20;
          13'h037B : pic_data = 24'hf10b0d;
          13'h037C : pic_data = 24'hf1180d;
          13'h037D : pic_data = 24'hf1230d;
          13'h037E : pic_data = 24'hf13b0d;
          13'h037F : pic_data = 24'hf1440d;
          13'h0380 : pic_data = 24'hf1520d;
          13'h0381 : pic_data = 24'hf15b0d;
          13'h0382 : pic_data = 24'hf1660d;
          13'h0383 : pic_data = 24'hf1800d;
          13'h0384 : pic_data = 24'hf1890d;
          13'h0385 : pic_data = 24'hf1970d;
          13'h0386 : pic_data = 24'hf1a00d;
          13'h0387 : pic_data = 24'hf1ab0d;
          13'h0388 : pic_data = 24'hf1c40d;
          13'h0389 : pic_data = 24'hf1cd0d;
          13'h038A : pic_data = 24'hf1db0d;
          13'h038B : pic_data = 24'hf1e40d;
          13'h038C : pic_data = 24'hf4f30d;
          13'h038D : pic_data = 24'hdbf10d;
          13'h038E : pic_data = 24'hd2f10d;
          13'h038F : pic_data = 24'hc5f10d;
          13'h0390 : pic_data = 24'hadf10d;
          13'h0391 : pic_data = 24'haef10d;
          13'h0392 : pic_data = 24'h99f10d;
          13'h0393 : pic_data = 24'h8ef10d;
          13'h0394 : pic_data = 24'h80f10d;
          13'h0395 : pic_data = 24'h68f10d;
          13'h0396 : pic_data = 24'h6af10d;
          13'h0397 : pic_data = 24'h54f10d;
          13'h0398 : pic_data = 24'h4af10d;
          13'h0399 : pic_data = 24'h3af10d;
          13'h039A : pic_data = 24'h25f10d;
          13'h039B : pic_data = 24'h26f10d;
          13'h039C : pic_data = 24'h0ff10c;
          13'h039D : pic_data = 24'h0cf113;
          13'h039E : pic_data = 24'h0df124;
          13'h039F : pic_data = 24'h0df137;
          13'h03A0 : pic_data = 24'h0df140;
          13'h03A1 : pic_data = 24'h0df153;
          13'h03A2 : pic_data = 24'h0df158;
          13'h03A3 : pic_data = 24'h0df167;
          13'h03A4 : pic_data = 24'h0df17b;
          13'h03A5 : pic_data = 24'h0df186;
          13'h03A6 : pic_data = 24'h0df198;
          13'h03A7 : pic_data = 24'h0df19b;
          13'h03A8 : pic_data = 24'h0df1ac;
          13'h03A9 : pic_data = 24'h0df1bf;
          13'h03AA : pic_data = 24'h0df1ca;
          13'h03AB : pic_data = 24'h0df1db;
          13'h03AC : pic_data = 24'h0df1df;
          13'h03AD : pic_data = 24'h0df3f3;
          13'h03AE : pic_data = 24'h0ddff1;
          13'h03AF : pic_data = 24'h0dd6f1;
          13'h03B0 : pic_data = 24'h0dc4f1;
          13'h03B1 : pic_data = 24'h0db2f1;
          13'h03B2 : pic_data = 24'h0dadf1;
          13'h03B3 : pic_data = 24'h0d9cf1;
          13'h03B4 : pic_data = 24'h0d92f1;
          13'h03B5 : pic_data = 24'h0d7ff1;
          13'h03B6 : pic_data = 24'h0d6df1;
          13'h03B7 : pic_data = 24'h0d69f1;
          13'h03B8 : pic_data = 24'h0d58f1;
          13'h03B9 : pic_data = 24'h0d4ff1;
          13'h03BA : pic_data = 24'h0d39f1;
          13'h03BB : pic_data = 24'h0d2af1;
          13'h03BC : pic_data = 24'h0d25f1;
          13'h03BD : pic_data = 24'h0c14f1;
          13'h03BE : pic_data = 24'h0f0cf1;
          13'h03BF : pic_data = 24'h240df1;
          13'h03C0 : pic_data = 24'h320df1;
          13'h03C1 : pic_data = 24'h3b0df1;
          13'h03C2 : pic_data = 24'h540df1;
          13'h03C3 : pic_data = 24'h530df1;
          13'h03C4 : pic_data = 24'h680df1;
          13'h03C5 : pic_data = 24'h770df1;
          13'h03C6 : pic_data = 24'h820df1;
          13'h03C7 : pic_data = 24'h990df1;
          13'h03C8 : pic_data = 24'h960df1;
          13'h03C9 : pic_data = 24'had0df1;
          13'h03CA : pic_data = 24'hbb0df1;
          13'h03CB : pic_data = 24'hc50df1;
          13'h03CC : pic_data = 24'hdc0df1;
          13'h03CD : pic_data = 24'hda0df1;
          13'h03CE : pic_data = 24'hf40df3;
          13'h03CF : pic_data = 24'hf10de4;
          13'h03D0 : pic_data = 24'hf10ddb;
          13'h03D1 : pic_data = 24'hf10dc3;
          13'h03D2 : pic_data = 24'hf10db7;
          13'h03D3 : pic_data = 24'hf10dac;
          13'h03D4 : pic_data = 24'hf10da0;
          13'h03D5 : pic_data = 24'hf10d97;
          13'h03D6 : pic_data = 24'hf10d7e;
          13'h03D7 : pic_data = 24'hf10d72;
          13'h03D8 : pic_data = 24'hf10d68;
          13'h03D9 : pic_data = 24'hf10d5b;
          13'h03DA : pic_data = 24'hf10d53;
          13'h03DB : pic_data = 24'hf10d38;
          13'h03DC : pic_data = 24'hf10d2f;
          13'h03DD : pic_data = 24'hf10d22;
          13'h03DE : pic_data = 24'hf20b0c;
          13'h03DF : pic_data = 24'hf2170c;
          13'h03E0 : pic_data = 24'hf2220c;
          13'h03E1 : pic_data = 24'hf23a0c;
          13'h03E2 : pic_data = 24'hf2440c;
          13'h03E3 : pic_data = 24'hf2520c;
          13'h03E4 : pic_data = 24'hf25b0c;
          13'h03E5 : pic_data = 24'hf2660c;
          13'h03E6 : pic_data = 24'hf2800c;
          13'h03E7 : pic_data = 24'hf2890c;
          13'h03E8 : pic_data = 24'hf2970c;
          13'h03E9 : pic_data = 24'hf2a00c;
          13'h03EA : pic_data = 24'hf2ab0c;
          13'h03EB : pic_data = 24'hf2c40c;
          13'h03EC : pic_data = 24'hf2ce0c;
          13'h03ED : pic_data = 24'hf2db0c;
          13'h03EE : pic_data = 24'hf2e50c;
          13'h03EF : pic_data = 24'hf5f40c;
          13'h03F0 : pic_data = 24'hdcf20c;
          13'h03F1 : pic_data = 24'hd2f20c;
          13'h03F2 : pic_data = 24'hc6f20c;
          13'h03F3 : pic_data = 24'hadf20c;
          13'h03F4 : pic_data = 24'haff20c;
          13'h03F5 : pic_data = 24'h99f20c;
          13'h03F6 : pic_data = 24'h8ef20c;
          13'h03F7 : pic_data = 24'h80f20c;
          13'h03F8 : pic_data = 24'h68f20c;
          13'h03F9 : pic_data = 24'h69f20c;
          13'h03FA : pic_data = 24'h53f20c;
          13'h03FB : pic_data = 24'h4af20c;
          13'h03FC : pic_data = 24'h39f20c;
          13'h03FD : pic_data = 24'h24f20c;
          13'h03FE : pic_data = 24'h25f20c;
          13'h03FF : pic_data = 24'h0ef20b;
          13'h0400 : pic_data = 24'h0cf212;
          13'h0401 : pic_data = 24'h0cf223;
          13'h0402 : pic_data = 24'h0cf236;
          13'h0403 : pic_data = 24'h0cf23f;
          13'h0404 : pic_data = 24'h0cf253;
          13'h0405 : pic_data = 24'h0cf257;
          13'h0406 : pic_data = 24'h0cf267;
          13'h0407 : pic_data = 24'h0cf27b;
          13'h0408 : pic_data = 24'h0cf286;
          13'h0409 : pic_data = 24'h0cf298;
          13'h040A : pic_data = 24'h0cf29b;
          13'h040B : pic_data = 24'h0cf2ac;
          13'h040C : pic_data = 24'h0cf2c0;
          13'h040D : pic_data = 24'h0cf2ca;
          13'h040E : pic_data = 24'h0cf2dc;
          13'h040F : pic_data = 24'h0cf2e0;
          13'h0410 : pic_data = 24'h0cf4f4;
          13'h0411 : pic_data = 24'h0ce0f2;
          13'h0412 : pic_data = 24'h0cd7f2;
          13'h0413 : pic_data = 24'h0cc5f2;
          13'h0414 : pic_data = 24'h0cb2f2;
          13'h0415 : pic_data = 24'h0caef2;
          13'h0416 : pic_data = 24'h0c9cf2;
          13'h0417 : pic_data = 24'h0c92f2;
          13'h0418 : pic_data = 24'h0c7ff2;
          13'h0419 : pic_data = 24'h0c6df2;
          13'h041A : pic_data = 24'h0c68f2;
          13'h041B : pic_data = 24'h0c58f2;
          13'h041C : pic_data = 24'h0c4ff2;
          13'h041D : pic_data = 24'h0c38f2;
          13'h041E : pic_data = 24'h0c29f2;
          13'h041F : pic_data = 24'h0c24f2;
          13'h0420 : pic_data = 24'h0c13f2;
          13'h0421 : pic_data = 24'h0e0bf2;
          13'h0422 : pic_data = 24'h240cf2;
          13'h0423 : pic_data = 24'h310cf2;
          13'h0424 : pic_data = 24'h3b0cf2;
          13'h0425 : pic_data = 24'h540cf2;
          13'h0426 : pic_data = 24'h520cf2;
          13'h0427 : pic_data = 24'h680cf2;
          13'h0428 : pic_data = 24'h770cf2;
          13'h0429 : pic_data = 24'h820cf2;
          13'h042A : pic_data = 24'h990cf2;
          13'h042B : pic_data = 24'h960cf2;
          13'h042C : pic_data = 24'had0cf2;
          13'h042D : pic_data = 24'hbb0cf2;
          13'h042E : pic_data = 24'hc60cf2;
          13'h042F : pic_data = 24'hdd0cf2;
          13'h0430 : pic_data = 24'hda0cf2;
          13'h0431 : pic_data = 24'hf50cf4;
          13'h0432 : pic_data = 24'hf20ce5;
          13'h0433 : pic_data = 24'hf20cdb;
          13'h0434 : pic_data = 24'hf20cc4;
          13'h0435 : pic_data = 24'hf20cb8;
          13'h0436 : pic_data = 24'hf20cad;
          13'h0437 : pic_data = 24'hf20ca0;
          13'h0438 : pic_data = 24'hf20c97;
          13'h0439 : pic_data = 24'hf20c7e;
          13'h043A : pic_data = 24'hf20c72;
          13'h043B : pic_data = 24'hf20c68;
          13'h043C : pic_data = 24'hf20c5b;
          13'h043D : pic_data = 24'hf20c53;
          13'h043E : pic_data = 24'hf20c37;
          13'h043F : pic_data = 24'hf20c2e;
          13'h0440 : pic_data = 24'hf20c22;
          13'h0441 : pic_data = 24'hed0f11;
          13'h0442 : pic_data = 24'hed1c11;
          13'h0443 : pic_data = 24'hed2511;
          13'h0444 : pic_data = 24'hed3f11;
          13'h0445 : pic_data = 24'hed4711;
          13'h0446 : pic_data = 24'hed5311;
          13'h0447 : pic_data = 24'hed5c11;
          13'h0448 : pic_data = 24'hed6711;
          13'h0449 : pic_data = 24'hed8011;
          13'h044A : pic_data = 24'hed8911;
          13'h044B : pic_data = 24'hed9611;
          13'h044C : pic_data = 24'hed9f11;
          13'h044D : pic_data = 24'hedaa11;
          13'h044E : pic_data = 24'hedc111;
          13'h044F : pic_data = 24'hedca11;
          13'h0450 : pic_data = 24'hedd811;
          13'h0451 : pic_data = 24'hede011;
          13'h0452 : pic_data = 24'hf0ef11;
          13'h0453 : pic_data = 24'hd8ed11;
          13'h0454 : pic_data = 24'hcfed11;
          13'h0455 : pic_data = 24'hc1ed11;
          13'h0456 : pic_data = 24'habed11;
          13'h0457 : pic_data = 24'haeed11;
          13'h0458 : pic_data = 24'h97ed11;
          13'h0459 : pic_data = 24'h8eed11;
          13'h045A : pic_data = 24'h80ed11;
          13'h045B : pic_data = 24'h69ed11;
          13'h045C : pic_data = 24'h6bed11;
          13'h045D : pic_data = 24'h54ed11;
          13'h045E : pic_data = 24'h4ced11;
          13'h045F : pic_data = 24'h3eed11;
          13'h0460 : pic_data = 24'h29ed11;
          13'h0461 : pic_data = 24'h28ed11;
          13'h0462 : pic_data = 24'h13ed10;
          13'h0463 : pic_data = 24'h10ed17;
          13'h0464 : pic_data = 24'h11ed26;
          13'h0465 : pic_data = 24'h11ed3b;
          13'h0466 : pic_data = 24'h11ed44;
          13'h0467 : pic_data = 24'h11ed53;
          13'h0468 : pic_data = 24'h11ed59;
          13'h0469 : pic_data = 24'h11ed68;
          13'h046A : pic_data = 24'h11ed7b;
          13'h046B : pic_data = 24'h11ed85;
          13'h046C : pic_data = 24'h11ed97;
          13'h046D : pic_data = 24'h11ed9a;
          13'h046E : pic_data = 24'h11edab;
          13'h046F : pic_data = 24'h11edbc;
          13'h0470 : pic_data = 24'h11edc6;
          13'h0471 : pic_data = 24'h11edd9;
          13'h0472 : pic_data = 24'h11eddb;
          13'h0473 : pic_data = 24'h11efef;
          13'h0474 : pic_data = 24'h11dded;
          13'h0475 : pic_data = 24'h11d3ed;
          13'h0476 : pic_data = 24'h11c0ed;
          13'h0477 : pic_data = 24'h11b0ed;
          13'h0478 : pic_data = 24'h11aded;
          13'h0479 : pic_data = 24'h119bed;
          13'h047A : pic_data = 24'h1191ed;
          13'h047B : pic_data = 24'h117fed;
          13'h047C : pic_data = 24'h116eed;
          13'h047D : pic_data = 24'h116aed;
          13'h047E : pic_data = 24'h1159ed;
          13'h047F : pic_data = 24'h114fed;
          13'h0480 : pic_data = 24'h113ded;
          13'h0481 : pic_data = 24'h112ced;
          13'h0482 : pic_data = 24'h1128ed;
          13'h0483 : pic_data = 24'h1017ed;
          13'h0484 : pic_data = 24'h1210ed;
          13'h0485 : pic_data = 24'h2711ed;
          13'h0486 : pic_data = 24'h3611ed;
          13'h0487 : pic_data = 24'h4011ed;
          13'h0488 : pic_data = 24'h5411ed;
          13'h0489 : pic_data = 24'h5411ed;
          13'h048A : pic_data = 24'h6911ed;
          13'h048B : pic_data = 24'h7711ed;
          13'h048C : pic_data = 24'h8211ed;
          13'h048D : pic_data = 24'h9811ed;
          13'h048E : pic_data = 24'h9511ed;
          13'h048F : pic_data = 24'hac11ed;
          13'h0490 : pic_data = 24'hb911ed;
          13'h0491 : pic_data = 24'hc111ed;
          13'h0492 : pic_data = 24'hda11ed;
          13'h0493 : pic_data = 24'hd711ed;
          13'h0494 : pic_data = 24'hf011ef;
          13'h0495 : pic_data = 24'hed11e0;
          13'h0496 : pic_data = 24'hed11d7;
          13'h0497 : pic_data = 24'hed11bf;
          13'h0498 : pic_data = 24'hed11b4;
          13'h0499 : pic_data = 24'hed11ac;
          13'h049A : pic_data = 24'hed119f;
          13'h049B : pic_data = 24'hed1196;
          13'h049C : pic_data = 24'hed117e;
          13'h049D : pic_data = 24'hed1173;
          13'h049E : pic_data = 24'hed1169;
          13'h049F : pic_data = 24'hed115c;
          13'h04A0 : pic_data = 24'hed1154;
          13'h04A1 : pic_data = 24'hed113c;
          13'h04A2 : pic_data = 24'hed1131;
          13'h04A3 : pic_data = 24'hed1125;
          13'h04A4 : pic_data = 24'hed0f11;
          13'h04A5 : pic_data = 24'hed1c11;
          13'h04A6 : pic_data = 24'hed2511;
          13'h04A7 : pic_data = 24'hed3f11;
          13'h04A8 : pic_data = 24'hed4711;
          13'h04A9 : pic_data = 24'hed5311;
          13'h04AA : pic_data = 24'hed5c11;
          13'h04AB : pic_data = 24'hed6711;
          13'h04AC : pic_data = 24'hed8011;
          13'h04AD : pic_data = 24'hed8911;
          13'h04AE : pic_data = 24'hed9611;
          13'h04AF : pic_data = 24'hed9f11;
          13'h04B0 : pic_data = 24'hedaa11;
          13'h04B1 : pic_data = 24'hedc111;
          13'h04B2 : pic_data = 24'hedca11;
          13'h04B3 : pic_data = 24'hedd811;
          13'h04B4 : pic_data = 24'hede011;
          13'h04B5 : pic_data = 24'hf0ef11;
          13'h04B6 : pic_data = 24'hd8ed11;
          13'h04B7 : pic_data = 24'hcfed11;
          13'h04B8 : pic_data = 24'hc1ed11;
          13'h04B9 : pic_data = 24'habed11;
          13'h04BA : pic_data = 24'haeed11;
          13'h04BB : pic_data = 24'h97ed11;
          13'h04BC : pic_data = 24'h8eed11;
          13'h04BD : pic_data = 24'h80ed11;
          13'h04BE : pic_data = 24'h69ed11;
          13'h04BF : pic_data = 24'h6bed11;
          13'h04C0 : pic_data = 24'h54ed11;
          13'h04C1 : pic_data = 24'h4ced11;
          13'h04C2 : pic_data = 24'h3eed11;
          13'h04C3 : pic_data = 24'h29ed11;
          13'h04C4 : pic_data = 24'h28ed11;
          13'h04C5 : pic_data = 24'h13ed10;
          13'h04C6 : pic_data = 24'h10ed17;
          13'h04C7 : pic_data = 24'h11ed26;
          13'h04C8 : pic_data = 24'h11ed3b;
          13'h04C9 : pic_data = 24'h11ed44;
          13'h04CA : pic_data = 24'h11ed53;
          13'h04CB : pic_data = 24'h11ed59;
          13'h04CC : pic_data = 24'h11ed68;
          13'h04CD : pic_data = 24'h11ed7b;
          13'h04CE : pic_data = 24'h11ed85;
          13'h04CF : pic_data = 24'h11ed97;
          13'h04D0 : pic_data = 24'h11ed9a;
          13'h04D1 : pic_data = 24'h11edab;
          13'h04D2 : pic_data = 24'h11edbc;
          13'h04D3 : pic_data = 24'h11edc6;
          13'h04D4 : pic_data = 24'h11edd9;
          13'h04D5 : pic_data = 24'h11eddb;
          13'h04D6 : pic_data = 24'h11eff0;
          13'h04D7 : pic_data = 24'h11dded;
          13'h04D8 : pic_data = 24'h11d3ed;
          13'h04D9 : pic_data = 24'h11c0ed;
          13'h04DA : pic_data = 24'h11b0ed;
          13'h04DB : pic_data = 24'h11aded;
          13'h04DC : pic_data = 24'h119bed;
          13'h04DD : pic_data = 24'h1191ed;
          13'h04DE : pic_data = 24'h117fed;
          13'h04DF : pic_data = 24'h116eed;
          13'h04E0 : pic_data = 24'h116aed;
          13'h04E1 : pic_data = 24'h1159ed;
          13'h04E2 : pic_data = 24'h114fed;
          13'h04E3 : pic_data = 24'h113ded;
          13'h04E4 : pic_data = 24'h112ced;
          13'h04E5 : pic_data = 24'h1128ed;
          13'h04E6 : pic_data = 24'h1017ed;
          13'h04E7 : pic_data = 24'h1210ed;
          13'h04E8 : pic_data = 24'h2711ed;
          13'h04E9 : pic_data = 24'h3611ed;
          13'h04EA : pic_data = 24'h4011ed;
          13'h04EB : pic_data = 24'h5411ed;
          13'h04EC : pic_data = 24'h5411ed;
          13'h04ED : pic_data = 24'h6911ed;
          13'h04EE : pic_data = 24'h7711ed;
          13'h04EF : pic_data = 24'h8211ed;
          13'h04F0 : pic_data = 24'h9811ed;
          13'h04F1 : pic_data = 24'h9511ed;
          13'h04F2 : pic_data = 24'hac11ed;
          13'h04F3 : pic_data = 24'hb911ed;
          13'h04F4 : pic_data = 24'hc111ed;
          13'h04F5 : pic_data = 24'hda11ed;
          13'h04F6 : pic_data = 24'hd711ed;
          13'h04F7 : pic_data = 24'hf011ef;
          13'h04F8 : pic_data = 24'hed11e0;
          13'h04F9 : pic_data = 24'hed11d7;
          13'h04FA : pic_data = 24'hed11bf;
          13'h04FB : pic_data = 24'hed11b4;
          13'h04FC : pic_data = 24'hed11ac;
          13'h04FD : pic_data = 24'hed119f;
          13'h04FE : pic_data = 24'hed1196;
          13'h04FF : pic_data = 24'hed117e;
          13'h0500 : pic_data = 24'hed1173;
          13'h0501 : pic_data = 24'hed1169;
          13'h0502 : pic_data = 24'hed115c;
          13'h0503 : pic_data = 24'hed1154;
          13'h0504 : pic_data = 24'hed113c;
          13'h0505 : pic_data = 24'hed1131;
          13'h0506 : pic_data = 24'hed1125;
          13'h0507 : pic_data = 24'hee0f10;
          13'h0508 : pic_data = 24'hee1b10;
          13'h0509 : pic_data = 24'hee2510;
          13'h050A : pic_data = 24'hee3f10;
          13'h050B : pic_data = 24'hee4710;
          13'h050C : pic_data = 24'hee5210;
          13'h050D : pic_data = 24'hee5c10;
          13'h050E : pic_data = 24'hee6710;
          13'h050F : pic_data = 24'hee8010;
          13'h0510 : pic_data = 24'hee8910;
          13'h0511 : pic_data = 24'hee9610;
          13'h0512 : pic_data = 24'hee9f10;
          13'h0513 : pic_data = 24'heeab10;
          13'h0514 : pic_data = 24'heec110;
          13'h0515 : pic_data = 24'heecb10;
          13'h0516 : pic_data = 24'heed810;
          13'h0517 : pic_data = 24'heee010;
          13'h0518 : pic_data = 24'hf0f010;
          13'h0519 : pic_data = 24'hd9ee10;
          13'h051A : pic_data = 24'hcfee10;
          13'h051B : pic_data = 24'hc1ee10;
          13'h051C : pic_data = 24'hacee10;
          13'h051D : pic_data = 24'haeee10;
          13'h051E : pic_data = 24'h98ee10;
          13'h051F : pic_data = 24'h8eee10;
          13'h0520 : pic_data = 24'h80ee10;
          13'h0521 : pic_data = 24'h69ee10;
          13'h0522 : pic_data = 24'h6aee10;
          13'h0523 : pic_data = 24'h54ee10;
          13'h0524 : pic_data = 24'h4cee10;
          13'h0525 : pic_data = 24'h3eee10;
          13'h0526 : pic_data = 24'h28ee10;
          13'h0527 : pic_data = 24'h28ee10;
          13'h0528 : pic_data = 24'h12ee0f;
          13'h0529 : pic_data = 24'h10ee16;
          13'h052A : pic_data = 24'h10ee26;
          13'h052B : pic_data = 24'h10ee3a;
          13'h052C : pic_data = 24'h10ee44;
          13'h052D : pic_data = 24'h10ee53;
          13'h052E : pic_data = 24'h10ee58;
          13'h052F : pic_data = 24'h10ee68;
          13'h0530 : pic_data = 24'h10ee7b;
          13'h0531 : pic_data = 24'h10ee85;
          13'h0532 : pic_data = 24'h10ee97;
          13'h0533 : pic_data = 24'h10ee9a;
          13'h0534 : pic_data = 24'h10eeac;
          13'h0535 : pic_data = 24'h10eebc;
          13'h0536 : pic_data = 24'h10eec6;
          13'h0537 : pic_data = 24'h10eed9;
          13'h0538 : pic_data = 24'h10eedb;
          13'h0539 : pic_data = 24'h10f0f0;
          13'h053A : pic_data = 24'h10ddee;
          13'h053B : pic_data = 24'h10d4ee;
          13'h053C : pic_data = 24'h10c0ee;
          13'h053D : pic_data = 24'h10b1ee;
          13'h053E : pic_data = 24'h10adee;
          13'h053F : pic_data = 24'h109bee;
          13'h0540 : pic_data = 24'h1091ee;
          13'h0541 : pic_data = 24'h107fee;
          13'h0542 : pic_data = 24'h106eee;
          13'h0543 : pic_data = 24'h1069ee;
          13'h0544 : pic_data = 24'h1059ee;
          13'h0545 : pic_data = 24'h104fee;
          13'h0546 : pic_data = 24'h103dee;
          13'h0547 : pic_data = 24'h102cee;
          13'h0548 : pic_data = 24'h1027ee;
          13'h0549 : pic_data = 24'h1016ee;
          13'h054A : pic_data = 24'h110fee;
          13'h054B : pic_data = 24'h2710ee;
          13'h054C : pic_data = 24'h3610ee;
          13'h054D : pic_data = 24'h3f10ee;
          13'h054E : pic_data = 24'h5410ee;
          13'h054F : pic_data = 24'h5310ee;
          13'h0550 : pic_data = 24'h6910ee;
          13'h0551 : pic_data = 24'h7710ee;
          13'h0552 : pic_data = 24'h8210ee;
          13'h0553 : pic_data = 24'h9810ee;
          13'h0554 : pic_data = 24'h9510ee;
          13'h0555 : pic_data = 24'had10ee;
          13'h0556 : pic_data = 24'hb910ee;
          13'h0557 : pic_data = 24'hc110ee;
          13'h0558 : pic_data = 24'hda10ee;
          13'h0559 : pic_data = 24'hd810ee;
          13'h055A : pic_data = 24'hf010f0;
          13'h055B : pic_data = 24'hee10e1;
          13'h055C : pic_data = 24'hee10d7;
          13'h055D : pic_data = 24'hee10c0;
          13'h055E : pic_data = 24'hee10b4;
          13'h055F : pic_data = 24'hee10ac;
          13'h0560 : pic_data = 24'hee10a0;
          13'h0561 : pic_data = 24'hee1096;
          13'h0562 : pic_data = 24'hee107e;
          13'h0563 : pic_data = 24'hee1073;
          13'h0564 : pic_data = 24'hee1069;
          13'h0565 : pic_data = 24'hee105c;
          13'h0566 : pic_data = 24'hee1054;
          13'h0567 : pic_data = 24'hee103c;
          13'h0568 : pic_data = 24'hee1031;
          13'h0569 : pic_data = 24'hee1025;
          13'h056A : pic_data = 24'he91315;
          13'h056B : pic_data = 24'he92015;
          13'h056C : pic_data = 24'he92915;
          13'h056D : pic_data = 24'he94115;
          13'h056E : pic_data = 24'he94915;
          13'h056F : pic_data = 24'he95515;
          13'h0570 : pic_data = 24'he95e15;
          13'h0571 : pic_data = 24'he96815;
          13'h0572 : pic_data = 24'he98015;
          13'h0573 : pic_data = 24'he98815;
          13'h0574 : pic_data = 24'he99515;
          13'h0575 : pic_data = 24'he99d15;
          13'h0576 : pic_data = 24'he9a815;
          13'h0577 : pic_data = 24'he9bf15;
          13'h0578 : pic_data = 24'he9c715;
          13'h0579 : pic_data = 24'he9d515;
          13'h057A : pic_data = 24'he9dd15;
          13'h057B : pic_data = 24'heceb15;
          13'h057C : pic_data = 24'hd5e915;
          13'h057D : pic_data = 24'hcce915;
          13'h057E : pic_data = 24'hbfe915;
          13'h057F : pic_data = 24'ha9e915;
          13'h0580 : pic_data = 24'hace915;
          13'h0581 : pic_data = 24'h95e915;
          13'h0582 : pic_data = 24'h8de915;
          13'h0583 : pic_data = 24'h80e915;
          13'h0584 : pic_data = 24'h6be915;
          13'h0585 : pic_data = 24'h6be915;
          13'h0586 : pic_data = 24'h57e915;
          13'h0587 : pic_data = 24'h4ee915;
          13'h0588 : pic_data = 24'h40e915;
          13'h0589 : pic_data = 24'h2ce915;
          13'h058A : pic_data = 24'h2ce915;
          13'h058B : pic_data = 24'h17e914;
          13'h058C : pic_data = 24'h14e91b;
          13'h058D : pic_data = 24'h15e92a;
          13'h058E : pic_data = 24'h15e93c;
          13'h058F : pic_data = 24'h15e946;
          13'h0590 : pic_data = 24'h15e956;
          13'h0591 : pic_data = 24'h15e959;
          13'h0592 : pic_data = 24'h15e969;
          13'h0593 : pic_data = 24'h15e97b;
          13'h0594 : pic_data = 24'h15e985;
          13'h0595 : pic_data = 24'h15e996;
          13'h0596 : pic_data = 24'h15e999;
          13'h0597 : pic_data = 24'h15e9a9;
          13'h0598 : pic_data = 24'h15e9ba;
          13'h0599 : pic_data = 24'h15e9c4;
          13'h059A : pic_data = 24'h15e9d6;
          13'h059B : pic_data = 24'h15e9d8;
          13'h059C : pic_data = 24'h15ebeb;
          13'h059D : pic_data = 24'h15d9e9;
          13'h059E : pic_data = 24'h15d0e9;
          13'h059F : pic_data = 24'h15bee9;
          13'h05A0 : pic_data = 24'h15aee9;
          13'h05A1 : pic_data = 24'h15abe9;
          13'h05A2 : pic_data = 24'h159ae9;
          13'h05A3 : pic_data = 24'h1591e9;
          13'h05A4 : pic_data = 24'h157fe9;
          13'h05A5 : pic_data = 24'h1570e9;
          13'h05A6 : pic_data = 24'h156ae9;
          13'h05A7 : pic_data = 24'h155be9;
          13'h05A8 : pic_data = 24'h1551e9;
          13'h05A9 : pic_data = 24'h153fe9;
          13'h05AA : pic_data = 24'h1531e9;
          13'h05AB : pic_data = 24'h152ce9;
          13'h05AC : pic_data = 24'h141be9;
          13'h05AD : pic_data = 24'h1614e9;
          13'h05AE : pic_data = 24'h2b15e9;
          13'h05AF : pic_data = 24'h3915e9;
          13'h05B0 : pic_data = 24'h4215e9;
          13'h05B1 : pic_data = 24'h5615e9;
          13'h05B2 : pic_data = 24'h5615e9;
          13'h05B3 : pic_data = 24'h6a15e9;
          13'h05B4 : pic_data = 24'h7815e9;
          13'h05B5 : pic_data = 24'h8015e9;
          13'h05B6 : pic_data = 24'h9715e9;
          13'h05B7 : pic_data = 24'h9415e9;
          13'h05B8 : pic_data = 24'haa15e9;
          13'h05B9 : pic_data = 24'hb715e9;
          13'h05BA : pic_data = 24'hbf15e9;
          13'h05BB : pic_data = 24'hd715e9;
          13'h05BC : pic_data = 24'hd415e9;
          13'h05BD : pic_data = 24'hec15eb;
          13'h05BE : pic_data = 24'he915dd;
          13'h05BF : pic_data = 24'he915d5;
          13'h05C0 : pic_data = 24'he915bd;
          13'h05C1 : pic_data = 24'he915b2;
          13'h05C2 : pic_data = 24'he915aa;
          13'h05C3 : pic_data = 24'he9159d;
          13'h05C4 : pic_data = 24'he91595;
          13'h05C5 : pic_data = 24'he9157e;
          13'h05C6 : pic_data = 24'he91573;
          13'h05C7 : pic_data = 24'he9156a;
          13'h05C8 : pic_data = 24'he9155e;
          13'h05C9 : pic_data = 24'he91556;
          13'h05CA : pic_data = 24'he9153e;
          13'h05CB : pic_data = 24'he91534;
          13'h05CC : pic_data = 24'he91529;
          13'h05CD : pic_data = 24'he91315;
          13'h05CE : pic_data = 24'he92015;
          13'h05CF : pic_data = 24'he92915;
          13'h05D0 : pic_data = 24'he94115;
          13'h05D1 : pic_data = 24'he94915;
          13'h05D2 : pic_data = 24'he95515;
          13'h05D3 : pic_data = 24'he95e15;
          13'h05D4 : pic_data = 24'he96815;
          13'h05D5 : pic_data = 24'he98015;
          13'h05D6 : pic_data = 24'he98815;
          13'h05D7 : pic_data = 24'he99515;
          13'h05D8 : pic_data = 24'he99d15;
          13'h05D9 : pic_data = 24'he9a815;
          13'h05DA : pic_data = 24'he9bf15;
          13'h05DB : pic_data = 24'he9c715;
          13'h05DC : pic_data = 24'he9d515;
          13'h05DD : pic_data = 24'he9dd15;
          13'h05DE : pic_data = 24'heceb15;
          13'h05DF : pic_data = 24'hd5e915;
          13'h05E0 : pic_data = 24'hcce915;
          13'h05E1 : pic_data = 24'hbfe915;
          13'h05E2 : pic_data = 24'ha9e915;
          13'h05E3 : pic_data = 24'hace915;
          13'h05E4 : pic_data = 24'h95e915;
          13'h05E5 : pic_data = 24'h8de915;
          13'h05E6 : pic_data = 24'h80e915;
          13'h05E7 : pic_data = 24'h6be915;
          13'h05E8 : pic_data = 24'h6be915;
          13'h05E9 : pic_data = 24'h57e915;
          13'h05EA : pic_data = 24'h4ee915;
          13'h05EB : pic_data = 24'h40e915;
          13'h05EC : pic_data = 24'h2ce915;
          13'h05ED : pic_data = 24'h2ce915;
          13'h05EE : pic_data = 24'h17e914;
          13'h05EF : pic_data = 24'h14e91b;
          13'h05F0 : pic_data = 24'h15e92a;
          13'h05F1 : pic_data = 24'h15e93c;
          13'h05F2 : pic_data = 24'h15e946;
          13'h05F3 : pic_data = 24'h15e956;
          13'h05F4 : pic_data = 24'h15e959;
          13'h05F5 : pic_data = 24'h15e969;
          13'h05F6 : pic_data = 24'h15e97b;
          13'h05F7 : pic_data = 24'h15e985;
          13'h05F8 : pic_data = 24'h15e996;
          13'h05F9 : pic_data = 24'h15e999;
          13'h05FA : pic_data = 24'h15e9a9;
          13'h05FB : pic_data = 24'h15e9ba;
          13'h05FC : pic_data = 24'h15e9c4;
          13'h05FD : pic_data = 24'h15e9d6;
          13'h05FE : pic_data = 24'h15e9d8;
          13'h05FF : pic_data = 24'h15ebeb;
          13'h0600 : pic_data = 24'h15d9e9;
          13'h0601 : pic_data = 24'h15d0e9;
          13'h0602 : pic_data = 24'h15bee9;
          13'h0603 : pic_data = 24'h15aee9;
          13'h0604 : pic_data = 24'h15abe9;
          13'h0605 : pic_data = 24'h159ae9;
          13'h0606 : pic_data = 24'h1591e9;
          13'h0607 : pic_data = 24'h157fe9;
          13'h0608 : pic_data = 24'h1570e9;
          13'h0609 : pic_data = 24'h156ae9;
          13'h060A : pic_data = 24'h155be9;
          13'h060B : pic_data = 24'h1551e9;
          13'h060C : pic_data = 24'h153fe9;
          13'h060D : pic_data = 24'h1531e9;
          13'h060E : pic_data = 24'h152ce9;
          13'h060F : pic_data = 24'h141be9;
          13'h0610 : pic_data = 24'h1614e9;
          13'h0611 : pic_data = 24'h2b15e9;
          13'h0612 : pic_data = 24'h3915e9;
          13'h0613 : pic_data = 24'h4215e9;
          13'h0614 : pic_data = 24'h5615e9;
          13'h0615 : pic_data = 24'h5615e9;
          13'h0616 : pic_data = 24'h6a15e9;
          13'h0617 : pic_data = 24'h7815e9;
          13'h0618 : pic_data = 24'h8015e9;
          13'h0619 : pic_data = 24'h9715e9;
          13'h061A : pic_data = 24'h9415e9;
          13'h061B : pic_data = 24'haa15e9;
          13'h061C : pic_data = 24'hb715e9;
          13'h061D : pic_data = 24'hbf15e9;
          13'h061E : pic_data = 24'hd715e9;
          13'h061F : pic_data = 24'hd415e9;
          13'h0620 : pic_data = 24'hec15eb;
          13'h0621 : pic_data = 24'he915dd;
          13'h0622 : pic_data = 24'he915d5;
          13'h0623 : pic_data = 24'he915bd;
          13'h0624 : pic_data = 24'he915b2;
          13'h0625 : pic_data = 24'he915aa;
          13'h0626 : pic_data = 24'he9159d;
          13'h0627 : pic_data = 24'he91595;
          13'h0628 : pic_data = 24'he9157f;
          13'h0629 : pic_data = 24'he91573;
          13'h062A : pic_data = 24'he9156a;
          13'h062B : pic_data = 24'he9155e;
          13'h062C : pic_data = 24'he91556;
          13'h062D : pic_data = 24'he9153e;
          13'h062E : pic_data = 24'he91534;
          13'h062F : pic_data = 24'he91529;
          13'h0630 : pic_data = 24'hea1314;
          13'h0631 : pic_data = 24'hea1f14;
          13'h0632 : pic_data = 24'hea2914;
          13'h0633 : pic_data = 24'hea4114;
          13'h0634 : pic_data = 24'hea4914;
          13'h0635 : pic_data = 24'hea5414;
          13'h0636 : pic_data = 24'hea5e14;
          13'h0637 : pic_data = 24'hea6814;
          13'h0638 : pic_data = 24'hea8014;
          13'h0639 : pic_data = 24'hea8814;
          13'h063A : pic_data = 24'hea9514;
          13'h063B : pic_data = 24'hea9d14;
          13'h063C : pic_data = 24'heaa914;
          13'h063D : pic_data = 24'heabf14;
          13'h063E : pic_data = 24'heac714;
          13'h063F : pic_data = 24'head514;
          13'h0640 : pic_data = 24'heade14;
          13'h0641 : pic_data = 24'heceb14;
          13'h0642 : pic_data = 24'hd6ea14;
          13'h0643 : pic_data = 24'hccea14;
          13'h0644 : pic_data = 24'hbfea14;
          13'h0645 : pic_data = 24'haaea14;
          13'h0646 : pic_data = 24'hacea14;
          13'h0647 : pic_data = 24'h95ea14;
          13'h0648 : pic_data = 24'h8dea14;
          13'h0649 : pic_data = 24'h80ea14;
          13'h064A : pic_data = 24'h6aea14;
          13'h064B : pic_data = 24'h6bea14;
          13'h064C : pic_data = 24'h56ea14;
          13'h064D : pic_data = 24'h4eea14;
          13'h064E : pic_data = 24'h40ea14;
          13'h064F : pic_data = 24'h2bea14;
          13'h0650 : pic_data = 24'h2cea14;
          13'h0651 : pic_data = 24'h16ea13;
          13'h0652 : pic_data = 24'h13ea1a;
          13'h0653 : pic_data = 24'h14ea2a;
          13'h0654 : pic_data = 24'h14ea3c;
          13'h0655 : pic_data = 24'h14ea46;
          13'h0656 : pic_data = 24'h14ea55;
          13'h0657 : pic_data = 24'h14ea59;
          13'h0658 : pic_data = 24'h14ea69;
          13'h0659 : pic_data = 24'h14ea7b;
          13'h065A : pic_data = 24'h14ea85;
          13'h065B : pic_data = 24'h14ea96;
          13'h065C : pic_data = 24'h14ea9a;
          13'h065D : pic_data = 24'h14eaaa;
          13'h065E : pic_data = 24'h14eaba;
          13'h065F : pic_data = 24'h14eac4;
          13'h0660 : pic_data = 24'h14ead6;
          13'h0661 : pic_data = 24'h14ead9;
          13'h0662 : pic_data = 24'h14ecec;
          13'h0663 : pic_data = 24'h14d9ea;
          13'h0664 : pic_data = 24'h14d1ea;
          13'h0665 : pic_data = 24'h14beea;
          13'h0666 : pic_data = 24'h14afea;
          13'h0667 : pic_data = 24'h14abea;
          13'h0668 : pic_data = 24'h149aea;
          13'h0669 : pic_data = 24'h1491ea;
          13'h066A : pic_data = 24'h147fea;
          13'h066B : pic_data = 24'h1470ea;
          13'h066C : pic_data = 24'h146aea;
          13'h066D : pic_data = 24'h145bea;
          13'h066E : pic_data = 24'h1451ea;
          13'h066F : pic_data = 24'h143fea;
          13'h0670 : pic_data = 24'h1430ea;
          13'h0671 : pic_data = 24'h142bea;
          13'h0672 : pic_data = 24'h141aea;
          13'h0673 : pic_data = 24'h1513ea;
          13'h0674 : pic_data = 24'h2b14ea;
          13'h0675 : pic_data = 24'h3914ea;
          13'h0676 : pic_data = 24'h4114ea;
          13'h0677 : pic_data = 24'h5614ea;
          13'h0678 : pic_data = 24'h5514ea;
          13'h0679 : pic_data = 24'h6a14ea;
          13'h067A : pic_data = 24'h7814ea;
          13'h067B : pic_data = 24'h8014ea;
          13'h067C : pic_data = 24'h9714ea;
          13'h067D : pic_data = 24'h9414ea;
          13'h067E : pic_data = 24'haa14ea;
          13'h067F : pic_data = 24'hb714ea;
          13'h0680 : pic_data = 24'hbf14ea;
          13'h0681 : pic_data = 24'hd714ea;
          13'h0682 : pic_data = 24'hd514ea;
          13'h0683 : pic_data = 24'hec14eb;
          13'h0684 : pic_data = 24'hea14de;
          13'h0685 : pic_data = 24'hea14d5;
          13'h0686 : pic_data = 24'hea14be;
          13'h0687 : pic_data = 24'hea14b2;
          13'h0688 : pic_data = 24'hea14aa;
          13'h0689 : pic_data = 24'hea149d;
          13'h068A : pic_data = 24'hea1495;
          13'h068B : pic_data = 24'hea147f;
          13'h068C : pic_data = 24'hea1473;
          13'h068D : pic_data = 24'hea146a;
          13'h068E : pic_data = 24'hea145e;
          13'h068F : pic_data = 24'hea1456;
          13'h0690 : pic_data = 24'hea143e;
          13'h0691 : pic_data = 24'hea1434;
          13'h0692 : pic_data = 24'hea1429;
          13'h0693 : pic_data = 24'he61819;
          13'h0694 : pic_data = 24'he62319;
          13'h0695 : pic_data = 24'he62c19;
          13'h0696 : pic_data = 24'he64319;
          13'h0697 : pic_data = 24'he64b19;
          13'h0698 : pic_data = 24'he65719;
          13'h0699 : pic_data = 24'he65f19;
          13'h069A : pic_data = 24'he66919;
          13'h069B : pic_data = 24'he68019;
          13'h069C : pic_data = 24'he68819;
          13'h069D : pic_data = 24'he69419;
          13'h069E : pic_data = 24'he69c19;
          13'h069F : pic_data = 24'he6a619;
          13'h06A0 : pic_data = 24'he6bd19;
          13'h06A1 : pic_data = 24'he6c519;
          13'h06A2 : pic_data = 24'he6d119;
          13'h06A3 : pic_data = 24'he6d919;
          13'h06A4 : pic_data = 24'he8e719;
          13'h06A5 : pic_data = 24'hd1e619;
          13'h06A6 : pic_data = 24'hc9e619;
          13'h06A7 : pic_data = 24'hbde619;
          13'h06A8 : pic_data = 24'ha7e619;
          13'h06A9 : pic_data = 24'haae619;
          13'h06AA : pic_data = 24'h94e619;
          13'h06AB : pic_data = 24'h8ce619;
          13'h06AC : pic_data = 24'h80e619;
          13'h06AD : pic_data = 24'h6ce619;
          13'h06AE : pic_data = 24'h6ce619;
          13'h06AF : pic_data = 24'h59e619;
          13'h06B0 : pic_data = 24'h50e619;
          13'h06B1 : pic_data = 24'h42e619;
          13'h06B2 : pic_data = 24'h2fe619;
          13'h06B3 : pic_data = 24'h2fe619;
          13'h06B4 : pic_data = 24'h1be619;
          13'h06B5 : pic_data = 24'h19e61e;
          13'h06B6 : pic_data = 24'h19e62d;
          13'h06B7 : pic_data = 24'h19e63e;
          13'h06B8 : pic_data = 24'h19e648;
          13'h06B9 : pic_data = 24'h19e657;
          13'h06BA : pic_data = 24'h19e65b;
          13'h06BB : pic_data = 24'h19e66a;
          13'h06BC : pic_data = 24'h19e67c;
          13'h06BD : pic_data = 24'h19e685;
          13'h06BE : pic_data = 24'h19e695;
          13'h06BF : pic_data = 24'h19e697;
          13'h06C0 : pic_data = 24'h19e6a7;
          13'h06C1 : pic_data = 24'h19e6b8;
          13'h06C2 : pic_data = 24'h19e6c1;
          13'h06C3 : pic_data = 24'h19e6d2;
          13'h06C4 : pic_data = 24'h19e6d4;
          13'h06C5 : pic_data = 24'h19e8e8;
          13'h06C6 : pic_data = 24'h19d5e6;
          13'h06C7 : pic_data = 24'h19cce6;
          13'h06C8 : pic_data = 24'h19bce6;
          13'h06C9 : pic_data = 24'h19ace6;
          13'h06CA : pic_data = 24'h19a9e6;
          13'h06CB : pic_data = 24'h1999e6;
          13'h06CC : pic_data = 24'h1990e6;
          13'h06CD : pic_data = 24'h197fe6;
          13'h06CE : pic_data = 24'h196fe6;
          13'h06CF : pic_data = 24'h196be6;
          13'h06D0 : pic_data = 24'h195ce6;
          13'h06D1 : pic_data = 24'h1953e6;
          13'h06D2 : pic_data = 24'h1941e6;
          13'h06D3 : pic_data = 24'h1932e6;
          13'h06D4 : pic_data = 24'h192ee6;
          13'h06D5 : pic_data = 24'h1920e6;
          13'h06D6 : pic_data = 24'h1b19e6;
          13'h06D7 : pic_data = 24'h2e19e6;
          13'h06D8 : pic_data = 24'h3b19e6;
          13'h06D9 : pic_data = 24'h4319e6;
          13'h06DA : pic_data = 24'h5819e6;
          13'h06DB : pic_data = 24'h5819e6;
          13'h06DC : pic_data = 24'h6b19e6;
          13'h06DD : pic_data = 24'h7819e6;
          13'h06DE : pic_data = 24'h8019e6;
          13'h06DF : pic_data = 24'h9619e6;
          13'h06E0 : pic_data = 24'h9319e6;
          13'h06E1 : pic_data = 24'ha819e6;
          13'h06E2 : pic_data = 24'hb519e6;
          13'h06E3 : pic_data = 24'hbd19e6;
          13'h06E4 : pic_data = 24'hd319e6;
          13'h06E5 : pic_data = 24'hd019e6;
          13'h06E6 : pic_data = 24'he819e7;
          13'h06E7 : pic_data = 24'he619d9;
          13'h06E8 : pic_data = 24'he619d1;
          13'h06E9 : pic_data = 24'he619bc;
          13'h06EA : pic_data = 24'he619b0;
          13'h06EB : pic_data = 24'he619a8;
          13'h06EC : pic_data = 24'he6199c;
          13'h06ED : pic_data = 24'he61994;
          13'h06EE : pic_data = 24'he6197f;
          13'h06EF : pic_data = 24'he61974;
          13'h06F0 : pic_data = 24'he6196b;
          13'h06F1 : pic_data = 24'he61960;
          13'h06F2 : pic_data = 24'he61958;
          13'h06F3 : pic_data = 24'he61940;
          13'h06F4 : pic_data = 24'he61937;
          13'h06F5 : pic_data = 24'he6192c;
          13'h06F6 : pic_data = 24'he5181a;
          13'h06F7 : pic_data = 24'he5241a;
          13'h06F8 : pic_data = 24'he52c1a;
          13'h06F9 : pic_data = 24'he5431a;
          13'h06FA : pic_data = 24'he54b1a;
          13'h06FB : pic_data = 24'he5571a;
          13'h06FC : pic_data = 24'he55f1a;
          13'h06FD : pic_data = 24'he5691a;
          13'h06FE : pic_data = 24'he5801a;
          13'h06FF : pic_data = 24'he5881a;
          13'h0700 : pic_data = 24'he5941a;
          13'h0701 : pic_data = 24'he59c1a;
          13'h0702 : pic_data = 24'he5a61a;
          13'h0703 : pic_data = 24'he5bd1a;
          13'h0704 : pic_data = 24'he5c51a;
          13'h0705 : pic_data = 24'he5d11a;
          13'h0706 : pic_data = 24'he5d91a;
          13'h0707 : pic_data = 24'he8e71a;
          13'h0708 : pic_data = 24'hd1e51a;
          13'h0709 : pic_data = 24'hc9e51a;
          13'h070A : pic_data = 24'hbde51a;
          13'h070B : pic_data = 24'ha7e51a;
          13'h070C : pic_data = 24'ha9e51a;
          13'h070D : pic_data = 24'h94e51a;
          13'h070E : pic_data = 24'h8ce51a;
          13'h070F : pic_data = 24'h80e51a;
          13'h0710 : pic_data = 24'h6ce51a;
          13'h0711 : pic_data = 24'h6ce51a;
          13'h0712 : pic_data = 24'h59e51a;
          13'h0713 : pic_data = 24'h50e51a;
          13'h0714 : pic_data = 24'h42e51a;
          13'h0715 : pic_data = 24'h2fe51a;
          13'h0716 : pic_data = 24'h2fe51a;
          13'h0717 : pic_data = 24'h1be519;
          13'h0718 : pic_data = 24'h19e51f;
          13'h0719 : pic_data = 24'h1ae52d;
          13'h071A : pic_data = 24'h1ae53e;
          13'h071B : pic_data = 24'h1ae548;
          13'h071C : pic_data = 24'h1ae558;
          13'h071D : pic_data = 24'h1ae55c;
          13'h071E : pic_data = 24'h1ae56a;
          13'h071F : pic_data = 24'h1ae57c;
          13'h0720 : pic_data = 24'h1ae585;
          13'h0721 : pic_data = 24'h1ae595;
          13'h0722 : pic_data = 24'h1ae597;
          13'h0723 : pic_data = 24'h1ae5a7;
          13'h0724 : pic_data = 24'h1ae5b8;
          13'h0725 : pic_data = 24'h1ae5c1;
          13'h0726 : pic_data = 24'h1ae5d2;
          13'h0727 : pic_data = 24'h1ae5d4;
          13'h0728 : pic_data = 24'h1ae7e7;
          13'h0729 : pic_data = 24'h1ad5e5;
          13'h072A : pic_data = 24'h1acce5;
          13'h072B : pic_data = 24'h1abce5;
          13'h072C : pic_data = 24'h1aace5;
          13'h072D : pic_data = 24'h1aa8e5;
          13'h072E : pic_data = 24'h1a99e5;
          13'h072F : pic_data = 24'h1a90e5;
          13'h0730 : pic_data = 24'h1a7fe5;
          13'h0731 : pic_data = 24'h1a6fe5;
          13'h0732 : pic_data = 24'h1a6ce5;
          13'h0733 : pic_data = 24'h1a5ce5;
          13'h0734 : pic_data = 24'h1a53e5;
          13'h0735 : pic_data = 24'h1a41e5;
          13'h0736 : pic_data = 24'h1a33e5;
          13'h0737 : pic_data = 24'h1a2ee5;
          13'h0738 : pic_data = 24'h1920e5;
          13'h0739 : pic_data = 24'h1b19e5;
          13'h073A : pic_data = 24'h2e1ae5;
          13'h073B : pic_data = 24'h3b1ae5;
          13'h073C : pic_data = 24'h441ae5;
          13'h073D : pic_data = 24'h581ae5;
          13'h073E : pic_data = 24'h581ae5;
          13'h073F : pic_data = 24'h6b1ae5;
          13'h0740 : pic_data = 24'h781ae5;
          13'h0741 : pic_data = 24'h811ae5;
          13'h0742 : pic_data = 24'h951ae5;
          13'h0743 : pic_data = 24'h931ae5;
          13'h0744 : pic_data = 24'ha81ae5;
          13'h0745 : pic_data = 24'hb51ae5;
          13'h0746 : pic_data = 24'hbd1ae5;
          13'h0747 : pic_data = 24'hd21ae5;
          13'h0748 : pic_data = 24'hd01ae5;
          13'h0749 : pic_data = 24'he81ae7;
          13'h074A : pic_data = 24'he51ad9;
          13'h074B : pic_data = 24'he51ad1;
          13'h074C : pic_data = 24'he51abc;
          13'h074D : pic_data = 24'he51ab0;
          13'h074E : pic_data = 24'he51aa8;
          13'h074F : pic_data = 24'he51a9c;
          13'h0750 : pic_data = 24'he51a94;
          13'h0751 : pic_data = 24'he51a7f;
          13'h0752 : pic_data = 24'he51a74;
          13'h0753 : pic_data = 24'he51a6b;
          13'h0754 : pic_data = 24'he51a61;
          13'h0755 : pic_data = 24'he51a58;
          13'h0756 : pic_data = 24'he51a40;
          13'h0757 : pic_data = 24'he51a38;
          13'h0758 : pic_data = 24'he51a2c;
          13'h0759 : pic_data = 24'he61819;
          13'h075A : pic_data = 24'he62319;
          13'h075B : pic_data = 24'he62c19;
          13'h075C : pic_data = 24'he64219;
          13'h075D : pic_data = 24'he64b19;
          13'h075E : pic_data = 24'he65719;
          13'h075F : pic_data = 24'he65f19;
          13'h0760 : pic_data = 24'he66919;
          13'h0761 : pic_data = 24'he68019;
          13'h0762 : pic_data = 24'he68819;
          13'h0763 : pic_data = 24'he69419;
          13'h0764 : pic_data = 24'he69c19;
          13'h0765 : pic_data = 24'he6a619;
          13'h0766 : pic_data = 24'he6bd19;
          13'h0767 : pic_data = 24'he6c619;
          13'h0768 : pic_data = 24'he6d119;
          13'h0769 : pic_data = 24'he6da19;
          13'h076A : pic_data = 24'he8e819;
          13'h076B : pic_data = 24'hd2e619;
          13'h076C : pic_data = 24'hc9e619;
          13'h076D : pic_data = 24'hbee619;
          13'h076E : pic_data = 24'ha7e619;
          13'h076F : pic_data = 24'haae619;
          13'h0770 : pic_data = 24'h95e619;
          13'h0771 : pic_data = 24'h8ce619;
          13'h0772 : pic_data = 24'h80e619;
          13'h0773 : pic_data = 24'h6ce619;
          13'h0774 : pic_data = 24'h6ce619;
          13'h0775 : pic_data = 24'h59e619;
          13'h0776 : pic_data = 24'h50e619;
          13'h0777 : pic_data = 24'h42e619;
          13'h0778 : pic_data = 24'h2ee619;
          13'h0779 : pic_data = 24'h2fe619;
          13'h077A : pic_data = 24'h1ae618;
          13'h077B : pic_data = 24'h19e61e;
          13'h077C : pic_data = 24'h19e62d;
          13'h077D : pic_data = 24'h19e63e;
          13'h077E : pic_data = 24'h19e648;
          13'h077F : pic_data = 24'h19e657;
          13'h0780 : pic_data = 24'h19e65b;
          13'h0781 : pic_data = 24'h19e66a;
          13'h0782 : pic_data = 24'h19e67c;
          13'h0783 : pic_data = 24'h19e685;
          13'h0784 : pic_data = 24'h19e695;
          13'h0785 : pic_data = 24'h19e697;
          13'h0786 : pic_data = 24'h19e6a7;
          13'h0787 : pic_data = 24'h19e6b8;
          13'h0788 : pic_data = 24'h19e6c1;
          13'h0789 : pic_data = 24'h19e6d2;
          13'h078A : pic_data = 24'h19e6d4;
          13'h078B : pic_data = 24'h19e8e8;
          13'h078C : pic_data = 24'h19d5e6;
          13'h078D : pic_data = 24'h19cce6;
          13'h078E : pic_data = 24'h19bde6;
          13'h078F : pic_data = 24'h19ade6;
          13'h0790 : pic_data = 24'h19a9e6;
          13'h0791 : pic_data = 24'h1999e6;
          13'h0792 : pic_data = 24'h1990e6;
          13'h0793 : pic_data = 24'h197fe6;
          13'h0794 : pic_data = 24'h196fe6;
          13'h0795 : pic_data = 24'h196be6;
          13'h0796 : pic_data = 24'h195ce6;
          13'h0797 : pic_data = 24'h1953e6;
          13'h0798 : pic_data = 24'h1941e6;
          13'h0799 : pic_data = 24'h1932e6;
          13'h079A : pic_data = 24'h192ee6;
          13'h079B : pic_data = 24'h191fe6;
          13'h079C : pic_data = 24'h1a18e6;
          13'h079D : pic_data = 24'h2e19e6;
          13'h079E : pic_data = 24'h3b19e6;
          13'h079F : pic_data = 24'h4319e6;
          13'h07A0 : pic_data = 24'h5819e6;
          13'h07A1 : pic_data = 24'h5819e6;
          13'h07A2 : pic_data = 24'h6b19e6;
          13'h07A3 : pic_data = 24'h7819e6;
          13'h07A4 : pic_data = 24'h8119e6;
          13'h07A5 : pic_data = 24'h9619e6;
          13'h07A6 : pic_data = 24'h9419e6;
          13'h07A7 : pic_data = 24'ha819e6;
          13'h07A8 : pic_data = 24'hb519e6;
          13'h07A9 : pic_data = 24'hbe19e6;
          13'h07AA : pic_data = 24'hd319e6;
          13'h07AB : pic_data = 24'hd119e6;
          13'h07AC : pic_data = 24'he819e8;
          13'h07AD : pic_data = 24'he619da;
          13'h07AE : pic_data = 24'he619d1;
          13'h07AF : pic_data = 24'he619bc;
          13'h07B0 : pic_data = 24'he619b0;
          13'h07B1 : pic_data = 24'he619a8;
          13'h07B2 : pic_data = 24'he6199c;
          13'h07B3 : pic_data = 24'he61994;
          13'h07B4 : pic_data = 24'he6197f;
          13'h07B5 : pic_data = 24'he61974;
          13'h07B6 : pic_data = 24'he6196a;
          13'h07B7 : pic_data = 24'he61960;
          13'h07B8 : pic_data = 24'he61958;
          13'h07B9 : pic_data = 24'he61940;
          13'h07BA : pic_data = 24'he61937;
          13'h07BB : pic_data = 24'he6192c;
          13'h07BC : pic_data = 24'he11c1d;
          13'h07BD : pic_data = 24'he1261d;
          13'h07BE : pic_data = 24'he12f1d;
          13'h07BF : pic_data = 24'he1461d;
          13'h07C0 : pic_data = 24'he14d1d;
          13'h07C1 : pic_data = 24'he1581d;
          13'h07C2 : pic_data = 24'he1601d;
          13'h07C3 : pic_data = 24'he16a1d;
          13'h07C4 : pic_data = 24'he1801d;
          13'h07C5 : pic_data = 24'he1881d;
          13'h07C6 : pic_data = 24'he1931d;
          13'h07C7 : pic_data = 24'he19b1d;
          13'h07C8 : pic_data = 24'he1a61d;
          13'h07C9 : pic_data = 24'he1ba1d;
          13'h07CA : pic_data = 24'he1c21d;
          13'h07CB : pic_data = 24'he1ce1d;
          13'h07CC : pic_data = 24'he1d51d;
          13'h07CD : pic_data = 24'he3e21d;
          13'h07CE : pic_data = 24'hcfe11d;
          13'h07CF : pic_data = 24'hc6e11d;
          13'h07D0 : pic_data = 24'hbae11d;
          13'h07D1 : pic_data = 24'ha7e11d;
          13'h07D2 : pic_data = 24'ha9e11d;
          13'h07D3 : pic_data = 24'h93e11d;
          13'h07D4 : pic_data = 24'h8ce11d;
          13'h07D5 : pic_data = 24'h80e11d;
          13'h07D6 : pic_data = 24'h6de11d;
          13'h07D7 : pic_data = 24'h6de11d;
          13'h07D8 : pic_data = 24'h5ae11d;
          13'h07D9 : pic_data = 24'h51e11d;
          13'h07DA : pic_data = 24'h45e11d;
          13'h07DB : pic_data = 24'h32e11d;
          13'h07DC : pic_data = 24'h32e11d;
          13'h07DD : pic_data = 24'h1fe11d;
          13'h07DE : pic_data = 24'h1de122;
          13'h07DF : pic_data = 24'h1de130;
          13'h07E0 : pic_data = 24'h1de141;
          13'h07E1 : pic_data = 24'h1de14a;
          13'h07E2 : pic_data = 24'h1de158;
          13'h07E3 : pic_data = 24'h1de15c;
          13'h07E4 : pic_data = 24'h1de16b;
          13'h07E5 : pic_data = 24'h1de17c;
          13'h07E6 : pic_data = 24'h1de184;
          13'h07E7 : pic_data = 24'h1de194;
          13'h07E8 : pic_data = 24'h1de196;
          13'h07E9 : pic_data = 24'h1de1a7;
          13'h07EA : pic_data = 24'h1de1b6;
          13'h07EB : pic_data = 24'h1de1be;
          13'h07EC : pic_data = 24'h1de1cf;
          13'h07ED : pic_data = 24'h1de1d1;
          13'h07EE : pic_data = 24'h1de2e2;
          13'h07EF : pic_data = 24'h1dd2e1;
          13'h07F0 : pic_data = 24'h1dc9e1;
          13'h07F1 : pic_data = 24'h1db9e1;
          13'h07F2 : pic_data = 24'h1daae1;
          13'h07F3 : pic_data = 24'h1da8e1;
          13'h07F4 : pic_data = 24'h1d98e1;
          13'h07F5 : pic_data = 24'h1d8fe1;
          13'h07F6 : pic_data = 24'h1d7fe1;
          13'h07F7 : pic_data = 24'h1d70e1;
          13'h07F8 : pic_data = 24'h1d6ce1;
          13'h07F9 : pic_data = 24'h1d5de1;
          13'h07FA : pic_data = 24'h1d55e1;
          13'h07FB : pic_data = 24'h1d44e1;
          13'h07FC : pic_data = 24'h1d35e1;
          13'h07FD : pic_data = 24'h1d31e1;
          13'h07FE : pic_data = 24'h1d23e1;
          13'h07FF : pic_data = 24'h1f1de1;
          13'h0800 : pic_data = 24'h311de1;
          13'h0801 : pic_data = 24'h3e1de1;
          13'h0802 : pic_data = 24'h471de1;
          13'h0803 : pic_data = 24'h591de1;
          13'h0804 : pic_data = 24'h591de1;
          13'h0805 : pic_data = 24'h6c1de1;
          13'h0806 : pic_data = 24'h781de1;
          13'h0807 : pic_data = 24'h811de1;
          13'h0808 : pic_data = 24'h941de1;
          13'h0809 : pic_data = 24'h931de1;
          13'h080A : pic_data = 24'ha71de1;
          13'h080B : pic_data = 24'hb21de1;
          13'h080C : pic_data = 24'hbb1de1;
          13'h080D : pic_data = 24'hd01de1;
          13'h080E : pic_data = 24'hce1de1;
          13'h080F : pic_data = 24'he31de2;
          13'h0810 : pic_data = 24'he11dd5;
          13'h0811 : pic_data = 24'he11dce;
          13'h0812 : pic_data = 24'he11db9;
          13'h0813 : pic_data = 24'he11dae;
          13'h0814 : pic_data = 24'he11da7;
          13'h0815 : pic_data = 24'he11d9b;
          13'h0816 : pic_data = 24'he11d93;
          13'h0817 : pic_data = 24'he11d7f;
          13'h0818 : pic_data = 24'he11d74;
          13'h0819 : pic_data = 24'he11d6c;
          13'h081A : pic_data = 24'he11d61;
          13'h081B : pic_data = 24'he11d59;
          13'h081C : pic_data = 24'he11d43;
          13'h081D : pic_data = 24'he11d3a;
          13'h081E : pic_data = 24'he11d2f;
          13'h081F : pic_data = 24'he11c1d;
          13'h0820 : pic_data = 24'he1261d;
          13'h0821 : pic_data = 24'he12f1d;
          13'h0822 : pic_data = 24'he1461d;
          13'h0823 : pic_data = 24'he14d1d;
          13'h0824 : pic_data = 24'he1581d;
          13'h0825 : pic_data = 24'he1601d;
          13'h0826 : pic_data = 24'he16b1d;
          13'h0827 : pic_data = 24'he1801d;
          13'h0828 : pic_data = 24'he1891d;
          13'h0829 : pic_data = 24'he1931d;
          13'h082A : pic_data = 24'he19b1d;
          13'h082B : pic_data = 24'he1a61d;
          13'h082C : pic_data = 24'he1ba1d;
          13'h082D : pic_data = 24'he1c21d;
          13'h082E : pic_data = 24'he1ce1d;
          13'h082F : pic_data = 24'he1d51d;
          13'h0830 : pic_data = 24'he3e21d;
          13'h0831 : pic_data = 24'hcfe11d;
          13'h0832 : pic_data = 24'hc6e11d;
          13'h0833 : pic_data = 24'hbae11d;
          13'h0834 : pic_data = 24'ha7e11d;
          13'h0835 : pic_data = 24'ha9e11d;
          13'h0836 : pic_data = 24'h93e11d;
          13'h0837 : pic_data = 24'h8ce11d;
          13'h0838 : pic_data = 24'h80e11d;
          13'h0839 : pic_data = 24'h6de11d;
          13'h083A : pic_data = 24'h6de11d;
          13'h083B : pic_data = 24'h5ae11d;
          13'h083C : pic_data = 24'h51e11d;
          13'h083D : pic_data = 24'h45e11d;
          13'h083E : pic_data = 24'h32e11d;
          13'h083F : pic_data = 24'h32e11d;
          13'h0840 : pic_data = 24'h1fe11d;
          13'h0841 : pic_data = 24'h1de123;
          13'h0842 : pic_data = 24'h1de130;
          13'h0843 : pic_data = 24'h1de141;
          13'h0844 : pic_data = 24'h1de14a;
          13'h0845 : pic_data = 24'h1de158;
          13'h0846 : pic_data = 24'h1de15c;
          13'h0847 : pic_data = 24'h1de16b;
          13'h0848 : pic_data = 24'h1de17c;
          13'h0849 : pic_data = 24'h1de184;
          13'h084A : pic_data = 24'h1de194;
          13'h084B : pic_data = 24'h1de196;
          13'h084C : pic_data = 24'h1de1a7;
          13'h084D : pic_data = 24'h1de1b6;
          13'h084E : pic_data = 24'h1de1be;
          13'h084F : pic_data = 24'h1de1cf;
          13'h0850 : pic_data = 24'h1de1d2;
          13'h0851 : pic_data = 24'h1de2e2;
          13'h0852 : pic_data = 24'h1dd2e1;
          13'h0853 : pic_data = 24'h1dc9e1;
          13'h0854 : pic_data = 24'h1db9e1;
          13'h0855 : pic_data = 24'h1daae1;
          13'h0856 : pic_data = 24'h1da8e1;
          13'h0857 : pic_data = 24'h1d98e1;
          13'h0858 : pic_data = 24'h1d8fe1;
          13'h0859 : pic_data = 24'h1d7fe1;
          13'h085A : pic_data = 24'h1d71e1;
          13'h085B : pic_data = 24'h1d6de1;
          13'h085C : pic_data = 24'h1d5de1;
          13'h085D : pic_data = 24'h1d55e1;
          13'h085E : pic_data = 24'h1d44e1;
          13'h085F : pic_data = 24'h1d35e1;
          13'h0860 : pic_data = 24'h1d31e1;
          13'h0861 : pic_data = 24'h1d22e1;
          13'h0862 : pic_data = 24'h1f1de1;
          13'h0863 : pic_data = 24'h311de1;
          13'h0864 : pic_data = 24'h3e1de1;
          13'h0865 : pic_data = 24'h471de1;
          13'h0866 : pic_data = 24'h591de1;
          13'h0867 : pic_data = 24'h591de1;
          13'h0868 : pic_data = 24'h6c1de1;
          13'h0869 : pic_data = 24'h781de1;
          13'h086A : pic_data = 24'h811de1;
          13'h086B : pic_data = 24'h941de1;
          13'h086C : pic_data = 24'h921de1;
          13'h086D : pic_data = 24'ha71de1;
          13'h086E : pic_data = 24'hb21de1;
          13'h086F : pic_data = 24'hbb1de1;
          13'h0870 : pic_data = 24'hd01de1;
          13'h0871 : pic_data = 24'hce1de1;
          13'h0872 : pic_data = 24'he31de2;
          13'h0873 : pic_data = 24'he11dd5;
          13'h0874 : pic_data = 24'he11dce;
          13'h0875 : pic_data = 24'he11db9;
          13'h0876 : pic_data = 24'he11dae;
          13'h0877 : pic_data = 24'he11da7;
          13'h0878 : pic_data = 24'he11d9b;
          13'h0879 : pic_data = 24'he11d92;
          13'h087A : pic_data = 24'he11d7f;
          13'h087B : pic_data = 24'he11d74;
          13'h087C : pic_data = 24'he11d6c;
          13'h087D : pic_data = 24'he11d61;
          13'h087E : pic_data = 24'he11d59;
          13'h087F : pic_data = 24'he11d43;
          13'h0880 : pic_data = 24'he11d3a;
          13'h0881 : pic_data = 24'he11d2f;
          13'h0882 : pic_data = 24'hdf1e1f;
          13'h0883 : pic_data = 24'hdf281f;
          13'h0884 : pic_data = 24'hdf311f;
          13'h0885 : pic_data = 24'hdf461f;
          13'h0886 : pic_data = 24'hdf4e1f;
          13'h0887 : pic_data = 24'hdf581f;
          13'h0888 : pic_data = 24'hdf611f;
          13'h0889 : pic_data = 24'hdf6a1f;
          13'h088A : pic_data = 24'hdf801f;
          13'h088B : pic_data = 24'hdf891f;
          13'h088C : pic_data = 24'hdf931f;
          13'h088D : pic_data = 24'hdf9b1f;
          13'h088E : pic_data = 24'hdfa51f;
          13'h088F : pic_data = 24'hdfb91f;
          13'h0890 : pic_data = 24'hdfc11f;
          13'h0891 : pic_data = 24'hdfcd1f;
          13'h0892 : pic_data = 24'hdfd41f;
          13'h0893 : pic_data = 24'he1e11f;
          13'h0894 : pic_data = 24'hcddf1f;
          13'h0895 : pic_data = 24'hc5df1f;
          13'h0896 : pic_data = 24'hbadf1f;
          13'h0897 : pic_data = 24'ha6df1f;
          13'h0898 : pic_data = 24'ha8df1f;
          13'h0899 : pic_data = 24'h93df1f;
          13'h089A : pic_data = 24'h8cdf1f;
          13'h089B : pic_data = 24'h80df1f;
          13'h089C : pic_data = 24'h6ddf1f;
          13'h089D : pic_data = 24'h6ddf1f;
          13'h089E : pic_data = 24'h5adf1f;
          13'h089F : pic_data = 24'h51df1f;
          13'h08A0 : pic_data = 24'h46df1f;
          13'h08A1 : pic_data = 24'h33df1f;
          13'h08A2 : pic_data = 24'h33df1f;
          13'h08A3 : pic_data = 24'h20df1e;
          13'h08A4 : pic_data = 24'h1edf24;
          13'h08A5 : pic_data = 24'h1fdf31;
          13'h08A6 : pic_data = 24'h1fdf42;
          13'h08A7 : pic_data = 24'h1fdf4b;
          13'h08A8 : pic_data = 24'h1fdf59;
          13'h08A9 : pic_data = 24'h1fdf5d;
          13'h08AA : pic_data = 24'h1fdf6b;
          13'h08AB : pic_data = 24'h1fdf7c;
          13'h08AC : pic_data = 24'h1fdf84;
          13'h08AD : pic_data = 24'h1fdf94;
          13'h08AE : pic_data = 24'h1fdf96;
          13'h08AF : pic_data = 24'h1fdfa6;
          13'h08B0 : pic_data = 24'h1fdfb6;
          13'h08B1 : pic_data = 24'h1fdfbd;
          13'h08B2 : pic_data = 24'h1fdfcd;
          13'h08B3 : pic_data = 24'h1fdfd0;
          13'h08B4 : pic_data = 24'h1fe1e1;
          13'h08B5 : pic_data = 24'h1fd1df;
          13'h08B6 : pic_data = 24'h1fc8df;
          13'h08B7 : pic_data = 24'h1fb9df;
          13'h08B8 : pic_data = 24'h1faadf;
          13'h08B9 : pic_data = 24'h1fa7df;
          13'h08BA : pic_data = 24'h1f98df;
          13'h08BB : pic_data = 24'h1f8fdf;
          13'h08BC : pic_data = 24'h1f7fdf;
          13'h08BD : pic_data = 24'h1f71df;
          13'h08BE : pic_data = 24'h1f6cdf;
          13'h08BF : pic_data = 24'h1f5edf;
          13'h08C0 : pic_data = 24'h1f56df;
          13'h08C1 : pic_data = 24'h1f45df;
          13'h08C2 : pic_data = 24'h1f37df;
          13'h08C3 : pic_data = 24'h1f33df;
          13'h08C4 : pic_data = 24'h1e24df;
          13'h08C5 : pic_data = 24'h201edf;
          13'h08C6 : pic_data = 24'h321fdf;
          13'h08C7 : pic_data = 24'h3f1fdf;
          13'h08C8 : pic_data = 24'h471fdf;
          13'h08C9 : pic_data = 24'h5a1fdf;
          13'h08CA : pic_data = 24'h591fdf;
          13'h08CB : pic_data = 24'h6c1fdf;
          13'h08CC : pic_data = 24'h781fdf;
          13'h08CD : pic_data = 24'h811fdf;
          13'h08CE : pic_data = 24'h941fdf;
          13'h08CF : pic_data = 24'h931fdf;
          13'h08D0 : pic_data = 24'ha71fdf;
          13'h08D1 : pic_data = 24'hb11fdf;
          13'h08D2 : pic_data = 24'hba1fdf;
          13'h08D3 : pic_data = 24'hce1fdf;
          13'h08D4 : pic_data = 24'hcc1fdf;
          13'h08D5 : pic_data = 24'he11fe1;
          13'h08D6 : pic_data = 24'hdf1fd4;
          13'h08D7 : pic_data = 24'hdf1fcc;
          13'h08D8 : pic_data = 24'hdf1fb8;
          13'h08D9 : pic_data = 24'hdf1fad;
          13'h08DA : pic_data = 24'hdf1fa6;
          13'h08DB : pic_data = 24'hdf1f9b;
          13'h08DC : pic_data = 24'hdf1f93;
          13'h08DD : pic_data = 24'hdf1f7f;
          13'h08DE : pic_data = 24'hdf1f74;
          13'h08DF : pic_data = 24'hdf1f6c;
          13'h08E0 : pic_data = 24'hdf1f62;
          13'h08E1 : pic_data = 24'hdf1f59;
          13'h08E2 : pic_data = 24'hdf1f44;
          13'h08E3 : pic_data = 24'hdf1f3b;
          13'h08E4 : pic_data = 24'hdf1f31;
          13'h08E5 : pic_data = 24'hdc2122;
          13'h08E6 : pic_data = 24'hdc2b22;
          13'h08E7 : pic_data = 24'hdc3422;
          13'h08E8 : pic_data = 24'hdc4822;
          13'h08E9 : pic_data = 24'hdc5022;
          13'h08EA : pic_data = 24'hdc5a22;
          13'h08EB : pic_data = 24'hdc6122;
          13'h08EC : pic_data = 24'hdc6a22;
          13'h08ED : pic_data = 24'hdc8022;
          13'h08EE : pic_data = 24'hdc8922;
          13'h08EF : pic_data = 24'hdc9322;
          13'h08F0 : pic_data = 24'hdc9a22;
          13'h08F1 : pic_data = 24'hdca322;
          13'h08F2 : pic_data = 24'hdcb722;
          13'h08F3 : pic_data = 24'hdcbf22;
          13'h08F4 : pic_data = 24'hdcc922;
          13'h08F5 : pic_data = 24'hdcd122;
          13'h08F6 : pic_data = 24'hdede22;
          13'h08F7 : pic_data = 24'hcadc22;
          13'h08F8 : pic_data = 24'hc3dc22;
          13'h08F9 : pic_data = 24'hb8dc22;
          13'h08FA : pic_data = 24'ha4dc22;
          13'h08FB : pic_data = 24'ha6dc22;
          13'h08FC : pic_data = 24'h94dc22;
          13'h08FD : pic_data = 24'h8cdc22;
          13'h08FE : pic_data = 24'h80dc22;
          13'h08FF : pic_data = 24'h6ddc22;
          13'h0900 : pic_data = 24'h6ddc22;
          13'h0901 : pic_data = 24'h5cdc22;
          13'h0902 : pic_data = 24'h53dc22;
          13'h0903 : pic_data = 24'h47dc22;
          13'h0904 : pic_data = 24'h36dc22;
          13'h0905 : pic_data = 24'h36dc22;
          13'h0906 : pic_data = 24'h23dc21;
          13'h0907 : pic_data = 24'h21dc27;
          13'h0908 : pic_data = 24'h22dc35;
          13'h0909 : pic_data = 24'h22dc44;
          13'h090A : pic_data = 24'h22dc4c;
          13'h090B : pic_data = 24'h22dc5b;
          13'h090C : pic_data = 24'h22dc5e;
          13'h090D : pic_data = 24'h22dc6b;
          13'h090E : pic_data = 24'h22dc7c;
          13'h090F : pic_data = 24'h22dc84;
          13'h0910 : pic_data = 24'h22dc94;
          13'h0911 : pic_data = 24'h22dc97;
          13'h0912 : pic_data = 24'h22dca4;
          13'h0913 : pic_data = 24'h22dcb4;
          13'h0914 : pic_data = 24'h22dcbc;
          13'h0915 : pic_data = 24'h22dcca;
          13'h0916 : pic_data = 24'h22dccd;
          13'h0917 : pic_data = 24'h22dede;
          13'h0918 : pic_data = 24'h22cedc;
          13'h0919 : pic_data = 24'h22c6dc;
          13'h091A : pic_data = 24'h22b7dc;
          13'h091B : pic_data = 24'h22a8dc;
          13'h091C : pic_data = 24'h22a5dc;
          13'h091D : pic_data = 24'h2297dc;
          13'h091E : pic_data = 24'h228fdc;
          13'h091F : pic_data = 24'h227fdc;
          13'h0920 : pic_data = 24'h2271dc;
          13'h0921 : pic_data = 24'h226cdc;
          13'h0922 : pic_data = 24'h225fdc;
          13'h0923 : pic_data = 24'h2258dc;
          13'h0924 : pic_data = 24'h2246dc;
          13'h0925 : pic_data = 24'h223adc;
          13'h0926 : pic_data = 24'h2236dc;
          13'h0927 : pic_data = 24'h2127dc;
          13'h0928 : pic_data = 24'h2321dc;
          13'h0929 : pic_data = 24'h3522dc;
          13'h092A : pic_data = 24'h4122dc;
          13'h092B : pic_data = 24'h4922dc;
          13'h092C : pic_data = 24'h5b22dc;
          13'h092D : pic_data = 24'h5a22dc;
          13'h092E : pic_data = 24'h6c22dc;
          13'h092F : pic_data = 24'h7822dc;
          13'h0930 : pic_data = 24'h8122dc;
          13'h0931 : pic_data = 24'h9422dc;
          13'h0932 : pic_data = 24'h9322dc;
          13'h0933 : pic_data = 24'ha522dc;
          13'h0934 : pic_data = 24'haf22dc;
          13'h0935 : pic_data = 24'hb922dc;
          13'h0936 : pic_data = 24'hcb22dc;
          13'h0937 : pic_data = 24'hc922dc;
          13'h0938 : pic_data = 24'hde22de;
          13'h0939 : pic_data = 24'hdc22d1;
          13'h093A : pic_data = 24'hdc22c9;
          13'h093B : pic_data = 24'hdc22b7;
          13'h093C : pic_data = 24'hdc22ac;
          13'h093D : pic_data = 24'hdc22a5;
          13'h093E : pic_data = 24'hdc229a;
          13'h093F : pic_data = 24'hdc2293;
          13'h0940 : pic_data = 24'hdc227f;
          13'h0941 : pic_data = 24'hdc2274;
          13'h0942 : pic_data = 24'hdc226c;
          13'h0943 : pic_data = 24'hdc2263;
          13'h0944 : pic_data = 24'hdc225b;
          13'h0945 : pic_data = 24'hdc2245;
          13'h0946 : pic_data = 24'hdc223e;
          13'h0947 : pic_data = 24'hdc2234;
          13'h0948 : pic_data = 24'hdd2021;
          13'h0949 : pic_data = 24'hdd2a21;
          13'h094A : pic_data = 24'hdd3321;
          13'h094B : pic_data = 24'hdd4721;
          13'h094C : pic_data = 24'hdd4f21;
          13'h094D : pic_data = 24'hdd5a21;
          13'h094E : pic_data = 24'hdd6121;
          13'h094F : pic_data = 24'hdd6a21;
          13'h0950 : pic_data = 24'hdd8021;
          13'h0951 : pic_data = 24'hdd8921;
          13'h0952 : pic_data = 24'hdd9321;
          13'h0953 : pic_data = 24'hdd9a21;
          13'h0954 : pic_data = 24'hdda421;
          13'h0955 : pic_data = 24'hddb821;
          13'h0956 : pic_data = 24'hddc021;
          13'h0957 : pic_data = 24'hddca21;
          13'h0958 : pic_data = 24'hddd121;
          13'h0959 : pic_data = 24'hdfde21;
          13'h095A : pic_data = 24'hcbdd21;
          13'h095B : pic_data = 24'hc3dd21;
          13'h095C : pic_data = 24'hb8dd21;
          13'h095D : pic_data = 24'ha5dd21;
          13'h095E : pic_data = 24'ha6dd21;
          13'h095F : pic_data = 24'h94dd21;
          13'h0960 : pic_data = 24'h8cdd21;
          13'h0961 : pic_data = 24'h80dd21;
          13'h0962 : pic_data = 24'h6ddd21;
          13'h0963 : pic_data = 24'h6ddd21;
          13'h0964 : pic_data = 24'h5cdd21;
          13'h0965 : pic_data = 24'h53dd21;
          13'h0966 : pic_data = 24'h47dd21;
          13'h0967 : pic_data = 24'h36dd21;
          13'h0968 : pic_data = 24'h36dd21;
          13'h0969 : pic_data = 24'h23dd21;
          13'h096A : pic_data = 24'h21dd26;
          13'h096B : pic_data = 24'h21dd34;
          13'h096C : pic_data = 24'h21dd44;
          13'h096D : pic_data = 24'h21dd4c;
          13'h096E : pic_data = 24'h21dd5a;
          13'h096F : pic_data = 24'h21dd5d;
          13'h0970 : pic_data = 24'h21dd6b;
          13'h0971 : pic_data = 24'h21dd7c;
          13'h0972 : pic_data = 24'h21dd84;
          13'h0973 : pic_data = 24'h21dd94;
          13'h0974 : pic_data = 24'h21dd97;
          13'h0975 : pic_data = 24'h21dda4;
          13'h0976 : pic_data = 24'h21ddb4;
          13'h0977 : pic_data = 24'h21ddbc;
          13'h0978 : pic_data = 24'h21ddcb;
          13'h0979 : pic_data = 24'h21ddce;
          13'h097A : pic_data = 24'h21dede;
          13'h097B : pic_data = 24'h21cedd;
          13'h097C : pic_data = 24'h21c6dd;
          13'h097D : pic_data = 24'h21b8dd;
          13'h097E : pic_data = 24'h21a8dd;
          13'h097F : pic_data = 24'h21a6dd;
          13'h0980 : pic_data = 24'h2197dd;
          13'h0981 : pic_data = 24'h218fdd;
          13'h0982 : pic_data = 24'h217fdd;
          13'h0983 : pic_data = 24'h2170dd;
          13'h0984 : pic_data = 24'h216cdd;
          13'h0985 : pic_data = 24'h215fdd;
          13'h0986 : pic_data = 24'h2157dd;
          13'h0987 : pic_data = 24'h2146dd;
          13'h0988 : pic_data = 24'h213add;
          13'h0989 : pic_data = 24'h2135dd;
          13'h098A : pic_data = 24'h2126dd;
          13'h098B : pic_data = 24'h2321dd;
          13'h098C : pic_data = 24'h3521dd;
          13'h098D : pic_data = 24'h4121dd;
          13'h098E : pic_data = 24'h4921dd;
          13'h098F : pic_data = 24'h5b21dd;
          13'h0990 : pic_data = 24'h5a21dd;
          13'h0991 : pic_data = 24'h6c21dd;
          13'h0992 : pic_data = 24'h7821dd;
          13'h0993 : pic_data = 24'h8121dd;
          13'h0994 : pic_data = 24'h9421dd;
          13'h0995 : pic_data = 24'h9321dd;
          13'h0996 : pic_data = 24'ha521dd;
          13'h0997 : pic_data = 24'hb021dd;
          13'h0998 : pic_data = 24'hb921dd;
          13'h0999 : pic_data = 24'hcb21dd;
          13'h099A : pic_data = 24'hca21dd;
          13'h099B : pic_data = 24'hdf21de;
          13'h099C : pic_data = 24'hdd21d1;
          13'h099D : pic_data = 24'hdd21ca;
          13'h099E : pic_data = 24'hdd21b7;
          13'h099F : pic_data = 24'hdd21ac;
          13'h09A0 : pic_data = 24'hdd21a5;
          13'h09A1 : pic_data = 24'hdd219a;
          13'h09A2 : pic_data = 24'hdd2193;
          13'h09A3 : pic_data = 24'hdd217f;
          13'h09A4 : pic_data = 24'hdd2174;
          13'h09A5 : pic_data = 24'hdd216b;
          13'h09A6 : pic_data = 24'hdd2162;
          13'h09A7 : pic_data = 24'hdd215b;
          13'h09A8 : pic_data = 24'hdd2145;
          13'h09A9 : pic_data = 24'hdd213d;
          13'h09AA : pic_data = 24'hdd2133;
          13'h09AB : pic_data = 24'hdb2223;
          13'h09AC : pic_data = 24'hdb2c23;
          13'h09AD : pic_data = 24'hdb3423;
          13'h09AE : pic_data = 24'hdb4923;
          13'h09AF : pic_data = 24'hdb5023;
          13'h09B0 : pic_data = 24'hdb5a23;
          13'h09B1 : pic_data = 24'hdb6223;
          13'h09B2 : pic_data = 24'hdb6b23;
          13'h09B3 : pic_data = 24'hdb8023;
          13'h09B4 : pic_data = 24'hdb8823;
          13'h09B5 : pic_data = 24'hdb9223;
          13'h09B6 : pic_data = 24'hdb9a23;
          13'h09B7 : pic_data = 24'hdba323;
          13'h09B8 : pic_data = 24'hdbb723;
          13'h09B9 : pic_data = 24'hdbbe23;
          13'h09BA : pic_data = 24'hdbc923;
          13'h09BB : pic_data = 24'hdbd023;
          13'h09BC : pic_data = 24'hdddd23;
          13'h09BD : pic_data = 24'hcadb23;
          13'h09BE : pic_data = 24'hc2db23;
          13'h09BF : pic_data = 24'hb7db23;
          13'h09C0 : pic_data = 24'ha4db23;
          13'h09C1 : pic_data = 24'ha6db23;
          13'h09C2 : pic_data = 24'h93db23;
          13'h09C3 : pic_data = 24'h8cdb23;
          13'h09C4 : pic_data = 24'h80db23;
          13'h09C5 : pic_data = 24'h6ddb23;
          13'h09C6 : pic_data = 24'h6ddb23;
          13'h09C7 : pic_data = 24'h5cdb23;
          13'h09C8 : pic_data = 24'h53db23;
          13'h09C9 : pic_data = 24'h48db23;
          13'h09CA : pic_data = 24'h37db23;
          13'h09CB : pic_data = 24'h37db23;
          13'h09CC : pic_data = 24'h24db22;
          13'h09CD : pic_data = 24'h22db28;
          13'h09CE : pic_data = 24'h23db35;
          13'h09CF : pic_data = 24'h23db45;
          13'h09D0 : pic_data = 24'h23db4d;
          13'h09D1 : pic_data = 24'h23db5b;
          13'h09D2 : pic_data = 24'h23db5e;
          13'h09D3 : pic_data = 24'h23db6b;
          13'h09D4 : pic_data = 24'h23db7c;
          13'h09D5 : pic_data = 24'h23db84;
          13'h09D6 : pic_data = 24'h23db93;
          13'h09D7 : pic_data = 24'h23db96;
          13'h09D8 : pic_data = 24'h23dba4;
          13'h09D9 : pic_data = 24'h23dbb3;
          13'h09DA : pic_data = 24'h23dbbb;
          13'h09DB : pic_data = 24'h23dbca;
          13'h09DC : pic_data = 24'h23dbcc;
          13'h09DD : pic_data = 24'h23dddd;
          13'h09DE : pic_data = 24'h23cddb;
          13'h09DF : pic_data = 24'h23c5db;
          13'h09E0 : pic_data = 24'h23b7db;
          13'h09E1 : pic_data = 24'h23a8db;
          13'h09E2 : pic_data = 24'h23a5db;
          13'h09E3 : pic_data = 24'h2397db;
          13'h09E4 : pic_data = 24'h238fdb;
          13'h09E5 : pic_data = 24'h237fdb;
          13'h09E6 : pic_data = 24'h2371db;
          13'h09E7 : pic_data = 24'h236ddb;
          13'h09E8 : pic_data = 24'h235fdb;
          13'h09E9 : pic_data = 24'h2358db;
          13'h09EA : pic_data = 24'h2347db;
          13'h09EB : pic_data = 24'h233bdb;
          13'h09EC : pic_data = 24'h2336db;
          13'h09ED : pic_data = 24'h2228db;
          13'h09EE : pic_data = 24'h2422db;
          13'h09EF : pic_data = 24'h3623db;
          13'h09F0 : pic_data = 24'h4223db;
          13'h09F1 : pic_data = 24'h4923db;
          13'h09F2 : pic_data = 24'h5c23db;
          13'h09F3 : pic_data = 24'h5a23db;
          13'h09F4 : pic_data = 24'h6c23db;
          13'h09F5 : pic_data = 24'h7823db;
          13'h09F6 : pic_data = 24'h8123db;
          13'h09F7 : pic_data = 24'h9423db;
          13'h09F8 : pic_data = 24'h9223db;
          13'h09F9 : pic_data = 24'ha523db;
          13'h09FA : pic_data = 24'haf23db;
          13'h09FB : pic_data = 24'hb823db;
          13'h09FC : pic_data = 24'hca23db;
          13'h09FD : pic_data = 24'hc823db;
          13'h09FE : pic_data = 24'hdd23dd;
          13'h09FF : pic_data = 24'hdb23d0;
          13'h0A00 : pic_data = 24'hdb23c9;
          13'h0A01 : pic_data = 24'hdb23b6;
          13'h0A02 : pic_data = 24'hdb23ac;
          13'h0A03 : pic_data = 24'hdb23a4;
          13'h0A04 : pic_data = 24'hdb239a;
          13'h0A05 : pic_data = 24'hdb2392;
          13'h0A06 : pic_data = 24'hdb237f;
          13'h0A07 : pic_data = 24'hdb2375;
          13'h0A08 : pic_data = 24'hdb236c;
          13'h0A09 : pic_data = 24'hdb2363;
          13'h0A0A : pic_data = 24'hdb235b;
          13'h0A0B : pic_data = 24'hdb2346;
          13'h0A0C : pic_data = 24'hdb233e;
          13'h0A0D : pic_data = 24'hdb2334;
          13'h0A0E : pic_data = 24'hd82526;
          13'h0A0F : pic_data = 24'hd82f26;
          13'h0A10 : pic_data = 24'hd83726;
          13'h0A11 : pic_data = 24'hd84b26;
          13'h0A12 : pic_data = 24'hd85226;
          13'h0A13 : pic_data = 24'hd85b26;
          13'h0A14 : pic_data = 24'hd86226;
          13'h0A15 : pic_data = 24'hd86c26;
          13'h0A16 : pic_data = 24'hd88026;
          13'h0A17 : pic_data = 24'hd88726;
          13'h0A18 : pic_data = 24'hd89226;
          13'h0A19 : pic_data = 24'hd89926;
          13'h0A1A : pic_data = 24'hd8a326;
          13'h0A1B : pic_data = 24'hd8b426;
          13'h0A1C : pic_data = 24'hd8bc26;
          13'h0A1D : pic_data = 24'hd8c726;
          13'h0A1E : pic_data = 24'hd8cd26;
          13'h0A1F : pic_data = 24'hdada26;
          13'h0A20 : pic_data = 24'hc7d826;
          13'h0A21 : pic_data = 24'hc0d826;
          13'h0A22 : pic_data = 24'hb5d826;
          13'h0A23 : pic_data = 24'ha4d826;
          13'h0A24 : pic_data = 24'ha5d826;
          13'h0A25 : pic_data = 24'h93d826;
          13'h0A26 : pic_data = 24'h8bd826;
          13'h0A27 : pic_data = 24'h80d826;
          13'h0A28 : pic_data = 24'h6ed826;
          13'h0A29 : pic_data = 24'h6ed826;
          13'h0A2A : pic_data = 24'h5dd826;
          13'h0A2B : pic_data = 24'h55d826;
          13'h0A2C : pic_data = 24'h4ad826;
          13'h0A2D : pic_data = 24'h39d826;
          13'h0A2E : pic_data = 24'h39d826;
          13'h0A2F : pic_data = 24'h27d825;
          13'h0A30 : pic_data = 24'h25d82b;
          13'h0A31 : pic_data = 24'h26d837;
          13'h0A32 : pic_data = 24'h26d848;
          13'h0A33 : pic_data = 24'h26d84e;
          13'h0A34 : pic_data = 24'h26d85b;
          13'h0A35 : pic_data = 24'h26d85f;
          13'h0A36 : pic_data = 24'h26d86c;
          13'h0A37 : pic_data = 24'h26d87c;
          13'h0A38 : pic_data = 24'h26d884;
          13'h0A39 : pic_data = 24'h26d892;
          13'h0A3A : pic_data = 24'h26d895;
          13'h0A3B : pic_data = 24'h26d8a3;
          13'h0A3C : pic_data = 24'h26d8b1;
          13'h0A3D : pic_data = 24'h26d8b9;
          13'h0A3E : pic_data = 24'h26d8c7;
          13'h0A3F : pic_data = 24'h26d8c9;
          13'h0A40 : pic_data = 24'h26dada;
          13'h0A41 : pic_data = 24'h26cbd8;
          13'h0A42 : pic_data = 24'h26c3d8;
          13'h0A43 : pic_data = 24'h26b4d8;
          13'h0A44 : pic_data = 24'h26a8d8;
          13'h0A45 : pic_data = 24'h26a4d8;
          13'h0A46 : pic_data = 24'h2696d8;
          13'h0A47 : pic_data = 24'h268ed8;
          13'h0A48 : pic_data = 24'h267fd8;
          13'h0A49 : pic_data = 24'h2672d8;
          13'h0A4A : pic_data = 24'h266dd8;
          13'h0A4B : pic_data = 24'h2660d8;
          13'h0A4C : pic_data = 24'h2658d8;
          13'h0A4D : pic_data = 24'h2649d8;
          13'h0A4E : pic_data = 24'h263dd8;
          13'h0A4F : pic_data = 24'h2638d8;
          13'h0A50 : pic_data = 24'h252bd8;
          13'h0A51 : pic_data = 24'h2725d8;
          13'h0A52 : pic_data = 24'h3826d8;
          13'h0A53 : pic_data = 24'h4426d8;
          13'h0A54 : pic_data = 24'h4b26d8;
          13'h0A55 : pic_data = 24'h5c26d8;
          13'h0A56 : pic_data = 24'h5b26d8;
          13'h0A57 : pic_data = 24'h6d26d8;
          13'h0A58 : pic_data = 24'h7926d8;
          13'h0A59 : pic_data = 24'h8126d8;
          13'h0A5A : pic_data = 24'h9326d8;
          13'h0A5B : pic_data = 24'h9226d8;
          13'h0A5C : pic_data = 24'ha426d8;
          13'h0A5D : pic_data = 24'had26d8;
          13'h0A5E : pic_data = 24'hb526d8;
          13'h0A5F : pic_data = 24'hc826d8;
          13'h0A60 : pic_data = 24'hc526d8;
          13'h0A61 : pic_data = 24'hda26d9;
          13'h0A62 : pic_data = 24'hd826ce;
          13'h0A63 : pic_data = 24'hd826c6;
          13'h0A64 : pic_data = 24'hd826b3;
          13'h0A65 : pic_data = 24'hd826ab;
          13'h0A66 : pic_data = 24'hd826a4;
          13'h0A67 : pic_data = 24'hd82699;
          13'h0A68 : pic_data = 24'hd82691;
          13'h0A69 : pic_data = 24'hd8267f;
          13'h0A6A : pic_data = 24'hd82675;
          13'h0A6B : pic_data = 24'hd8266d;
          13'h0A6C : pic_data = 24'hd82664;
          13'h0A6D : pic_data = 24'hd8265c;
          13'h0A6E : pic_data = 24'hd82649;
          13'h0A6F : pic_data = 24'hd82641;
          13'h0A70 : pic_data = 24'hd82637;
          13'h0A71 : pic_data = 24'hd92425;
          13'h0A72 : pic_data = 24'hd92e25;
          13'h0A73 : pic_data = 24'hd93625;
          13'h0A74 : pic_data = 24'hd94b25;
          13'h0A75 : pic_data = 24'hd95125;
          13'h0A76 : pic_data = 24'hd95b25;
          13'h0A77 : pic_data = 24'hd96225;
          13'h0A78 : pic_data = 24'hd96b25;
          13'h0A79 : pic_data = 24'hd98025;
          13'h0A7A : pic_data = 24'hd98725;
          13'h0A7B : pic_data = 24'hd99225;
          13'h0A7C : pic_data = 24'hd99925;
          13'h0A7D : pic_data = 24'hd9a325;
          13'h0A7E : pic_data = 24'hd9b425;
          13'h0A7F : pic_data = 24'hd9bc25;
          13'h0A80 : pic_data = 24'hd9c725;
          13'h0A81 : pic_data = 24'hd9cd25;
          13'h0A82 : pic_data = 24'hdbda25;
          13'h0A83 : pic_data = 24'hc8d925;
          13'h0A84 : pic_data = 24'hc0d925;
          13'h0A85 : pic_data = 24'hb5d925;
          13'h0A86 : pic_data = 24'ha4d925;
          13'h0A87 : pic_data = 24'ha5d925;
          13'h0A88 : pic_data = 24'h93d925;
          13'h0A89 : pic_data = 24'h8bd925;
          13'h0A8A : pic_data = 24'h80d925;
          13'h0A8B : pic_data = 24'h6ed925;
          13'h0A8C : pic_data = 24'h6ed925;
          13'h0A8D : pic_data = 24'h5dd925;
          13'h0A8E : pic_data = 24'h55d925;
          13'h0A8F : pic_data = 24'h4ad925;
          13'h0A90 : pic_data = 24'h39d925;
          13'h0A91 : pic_data = 24'h39d925;
          13'h0A92 : pic_data = 24'h27d925;
          13'h0A93 : pic_data = 24'h25d92b;
          13'h0A94 : pic_data = 24'h25d937;
          13'h0A95 : pic_data = 24'h25d947;
          13'h0A96 : pic_data = 24'h25d94e;
          13'h0A97 : pic_data = 24'h25d95b;
          13'h0A98 : pic_data = 24'h25d95e;
          13'h0A99 : pic_data = 24'h25d96c;
          13'h0A9A : pic_data = 24'h25d97c;
          13'h0A9B : pic_data = 24'h25d984;
          13'h0A9C : pic_data = 24'h25d993;
          13'h0A9D : pic_data = 24'h25d996;
          13'h0A9E : pic_data = 24'h25d9a4;
          13'h0A9F : pic_data = 24'h25d9b1;
          13'h0AA0 : pic_data = 24'h25d9b9;
          13'h0AA1 : pic_data = 24'h25d9c8;
          13'h0AA2 : pic_data = 24'h25d9c9;
          13'h0AA3 : pic_data = 24'h25dada;
          13'h0AA4 : pic_data = 24'h25cbd9;
          13'h0AA5 : pic_data = 24'h25c3d9;
          13'h0AA6 : pic_data = 24'h25b4d9;
          13'h0AA7 : pic_data = 24'h25a8d9;
          13'h0AA8 : pic_data = 24'h25a5d9;
          13'h0AA9 : pic_data = 24'h2596d9;
          13'h0AAA : pic_data = 24'h258ed9;
          13'h0AAB : pic_data = 24'h257fd9;
          13'h0AAC : pic_data = 24'h2572d9;
          13'h0AAD : pic_data = 24'h256dd9;
          13'h0AAE : pic_data = 24'h2560d9;
          13'h0AAF : pic_data = 24'h2558d9;
          13'h0AB0 : pic_data = 24'h2549d9;
          13'h0AB1 : pic_data = 24'h253dd9;
          13'h0AB2 : pic_data = 24'h2538d9;
          13'h0AB3 : pic_data = 24'h252bd9;
          13'h0AB4 : pic_data = 24'h2725d9;
          13'h0AB5 : pic_data = 24'h3825d9;
          13'h0AB6 : pic_data = 24'h4425d9;
          13'h0AB7 : pic_data = 24'h4b25d9;
          13'h0AB8 : pic_data = 24'h5c25d9;
          13'h0AB9 : pic_data = 24'h5b25d9;
          13'h0ABA : pic_data = 24'h6d25d9;
          13'h0ABB : pic_data = 24'h7925d9;
          13'h0ABC : pic_data = 24'h8125d9;
          13'h0ABD : pic_data = 24'h9325d9;
          13'h0ABE : pic_data = 24'h9225d9;
          13'h0ABF : pic_data = 24'ha425d9;
          13'h0AC0 : pic_data = 24'hae25d9;
          13'h0AC1 : pic_data = 24'hb625d9;
          13'h0AC2 : pic_data = 24'hc825d9;
          13'h0AC3 : pic_data = 24'hc625d9;
          13'h0AC4 : pic_data = 24'hdb25da;
          13'h0AC5 : pic_data = 24'hd925cf;
          13'h0AC6 : pic_data = 24'hd925c7;
          13'h0AC7 : pic_data = 24'hd925b4;
          13'h0AC8 : pic_data = 24'hd925ab;
          13'h0AC9 : pic_data = 24'hd925a4;
          13'h0ACA : pic_data = 24'hd92599;
          13'h0ACB : pic_data = 24'hd92592;
          13'h0ACC : pic_data = 24'hd9257f;
          13'h0ACD : pic_data = 24'hd92575;
          13'h0ACE : pic_data = 24'hd9256c;
          13'h0ACF : pic_data = 24'hd92563;
          13'h0AD0 : pic_data = 24'hd9255b;
          13'h0AD1 : pic_data = 24'hd92548;
          13'h0AD2 : pic_data = 24'hd92540;
          13'h0AD3 : pic_data = 24'hd92536;
          13'h0AD4 : pic_data = 24'hd72627;
          13'h0AD5 : pic_data = 24'hd73027;
          13'h0AD6 : pic_data = 24'hd73827;
          13'h0AD7 : pic_data = 24'hd74c27;
          13'h0AD8 : pic_data = 24'hd75227;
          13'h0AD9 : pic_data = 24'hd75b27;
          13'h0ADA : pic_data = 24'hd76327;
          13'h0ADB : pic_data = 24'hd76c27;
          13'h0ADC : pic_data = 24'hd78027;
          13'h0ADD : pic_data = 24'hd78727;
          13'h0ADE : pic_data = 24'hd79127;
          13'h0ADF : pic_data = 24'hd79927;
          13'h0AE0 : pic_data = 24'hd7a227;
          13'h0AE1 : pic_data = 24'hd7b427;
          13'h0AE2 : pic_data = 24'hd7bc27;
          13'h0AE3 : pic_data = 24'hd7c627;
          13'h0AE4 : pic_data = 24'hd7cc27;
          13'h0AE5 : pic_data = 24'hd9d927;
          13'h0AE6 : pic_data = 24'hc7d727;
          13'h0AE7 : pic_data = 24'hbfd727;
          13'h0AE8 : pic_data = 24'hb4d727;
          13'h0AE9 : pic_data = 24'ha3d727;
          13'h0AEA : pic_data = 24'ha5d727;
          13'h0AEB : pic_data = 24'h92d727;
          13'h0AEC : pic_data = 24'h8bd727;
          13'h0AED : pic_data = 24'h80d727;
          13'h0AEE : pic_data = 24'h6ed727;
          13'h0AEF : pic_data = 24'h6fd727;
          13'h0AF0 : pic_data = 24'h5dd727;
          13'h0AF1 : pic_data = 24'h56d727;
          13'h0AF2 : pic_data = 24'h4bd727;
          13'h0AF3 : pic_data = 24'h3ad727;
          13'h0AF4 : pic_data = 24'h3ad727;
          13'h0AF5 : pic_data = 24'h28d726;
          13'h0AF6 : pic_data = 24'h27d72c;
          13'h0AF7 : pic_data = 24'h27d738;
          13'h0AF8 : pic_data = 24'h27d748;
          13'h0AF9 : pic_data = 24'h27d74f;
          13'h0AFA : pic_data = 24'h27d75c;
          13'h0AFB : pic_data = 24'h27d75f;
          13'h0AFC : pic_data = 24'h27d76d;
          13'h0AFD : pic_data = 24'h27d77c;
          13'h0AFE : pic_data = 24'h27d784;
          13'h0AFF : pic_data = 24'h27d792;
          13'h0B00 : pic_data = 24'h27d795;
          13'h0B01 : pic_data = 24'h27d7a3;
          13'h0B02 : pic_data = 24'h27d7b0;
          13'h0B03 : pic_data = 24'h27d7b8;
          13'h0B04 : pic_data = 24'h27d7c7;
          13'h0B05 : pic_data = 24'h27d7c8;
          13'h0B06 : pic_data = 24'h27d9d9;
          13'h0B07 : pic_data = 24'h27cad7;
          13'h0B08 : pic_data = 24'h27c2d7;
          13'h0B09 : pic_data = 24'h27b4d7;
          13'h0B0A : pic_data = 24'h27a7d7;
          13'h0B0B : pic_data = 24'h27a4d7;
          13'h0B0C : pic_data = 24'h2796d7;
          13'h0B0D : pic_data = 24'h278ed7;
          13'h0B0E : pic_data = 24'h277fd7;
          13'h0B0F : pic_data = 24'h2772d7;
          13'h0B10 : pic_data = 24'h276ed7;
          13'h0B11 : pic_data = 24'h2761d7;
          13'h0B12 : pic_data = 24'h2759d7;
          13'h0B13 : pic_data = 24'h274ad7;
          13'h0B14 : pic_data = 24'h273ed7;
          13'h0B15 : pic_data = 24'h2739d7;
          13'h0B16 : pic_data = 24'h272cd7;
          13'h0B17 : pic_data = 24'h2826d7;
          13'h0B18 : pic_data = 24'h3927d7;
          13'h0B19 : pic_data = 24'h4527d7;
          13'h0B1A : pic_data = 24'h4b27d7;
          13'h0B1B : pic_data = 24'h5d27d7;
          13'h0B1C : pic_data = 24'h5c27d7;
          13'h0B1D : pic_data = 24'h6e27d7;
          13'h0B1E : pic_data = 24'h7927d7;
          13'h0B1F : pic_data = 24'h8127d7;
          13'h0B20 : pic_data = 24'h9327d7;
          13'h0B21 : pic_data = 24'h9227d7;
          13'h0B22 : pic_data = 24'ha427d7;
          13'h0B23 : pic_data = 24'had27d7;
          13'h0B24 : pic_data = 24'hb527d7;
          13'h0B25 : pic_data = 24'hc827d7;
          13'h0B26 : pic_data = 24'hc527d7;
          13'h0B27 : pic_data = 24'hd927d9;
          13'h0B28 : pic_data = 24'hd727cd;
          13'h0B29 : pic_data = 24'hd727c6;
          13'h0B2A : pic_data = 24'hd727b3;
          13'h0B2B : pic_data = 24'hd727ab;
          13'h0B2C : pic_data = 24'hd727a3;
          13'h0B2D : pic_data = 24'hd72799;
          13'h0B2E : pic_data = 24'hd72791;
          13'h0B2F : pic_data = 24'hd7277f;
          13'h0B30 : pic_data = 24'hd72776;
          13'h0B31 : pic_data = 24'hd7276d;
          13'h0B32 : pic_data = 24'hd72764;
          13'h0B33 : pic_data = 24'hd7275c;
          13'h0B34 : pic_data = 24'hd72749;
          13'h0B35 : pic_data = 24'hd72741;
          13'h0B36 : pic_data = 24'hd72738;
          13'h0B37 : pic_data = 24'hd42a2b;
          13'h0B38 : pic_data = 24'hd4332b;
          13'h0B39 : pic_data = 24'hd43b2b;
          13'h0B3A : pic_data = 24'hd44e2b;
          13'h0B3B : pic_data = 24'hd4552b;
          13'h0B3C : pic_data = 24'hd45e2b;
          13'h0B3D : pic_data = 24'hd4662b;
          13'h0B3E : pic_data = 24'hd46e2b;
          13'h0B3F : pic_data = 24'hd47f2b;
          13'h0B40 : pic_data = 24'hd4882b;
          13'h0B41 : pic_data = 24'hd4912b;
          13'h0B42 : pic_data = 24'hd4982b;
          13'h0B43 : pic_data = 24'hd4a02b;
          13'h0B44 : pic_data = 24'hd4b22b;
          13'h0B45 : pic_data = 24'hd4b92b;
          13'h0B46 : pic_data = 24'hd4c42b;
          13'h0B47 : pic_data = 24'hd4ca2b;
          13'h0B48 : pic_data = 24'hd6d52b;
          13'h0B49 : pic_data = 24'hc4d42b;
          13'h0B4A : pic_data = 24'hbcd42b;
          13'h0B4B : pic_data = 24'hb3d42b;
          13'h0B4C : pic_data = 24'ha2d42b;
          13'h0B4D : pic_data = 24'ha3d42b;
          13'h0B4E : pic_data = 24'h92d42b;
          13'h0B4F : pic_data = 24'h8bd42b;
          13'h0B50 : pic_data = 24'h80d42b;
          13'h0B51 : pic_data = 24'h6fd42b;
          13'h0B52 : pic_data = 24'h70d42b;
          13'h0B53 : pic_data = 24'h5fd42b;
          13'h0B54 : pic_data = 24'h58d42b;
          13'h0B55 : pic_data = 24'h4dd42b;
          13'h0B56 : pic_data = 24'h3dd42b;
          13'h0B57 : pic_data = 24'h3dd42b;
          13'h0B58 : pic_data = 24'h2dd42a;
          13'h0B59 : pic_data = 24'h2bd430;
          13'h0B5A : pic_data = 24'h2bd43b;
          13'h0B5B : pic_data = 24'h2bd44b;
          13'h0B5C : pic_data = 24'h2bd451;
          13'h0B5D : pic_data = 24'h2bd45f;
          13'h0B5E : pic_data = 24'h2bd462;
          13'h0B5F : pic_data = 24'h2bd46f;
          13'h0B60 : pic_data = 24'h2bd47c;
          13'h0B61 : pic_data = 24'h2bd484;
          13'h0B62 : pic_data = 24'h2bd491;
          13'h0B63 : pic_data = 24'h2bd495;
          13'h0B64 : pic_data = 24'h2bd4a1;
          13'h0B65 : pic_data = 24'h2bd4af;
          13'h0B66 : pic_data = 24'h2bd4b6;
          13'h0B67 : pic_data = 24'h2bd4c4;
          13'h0B68 : pic_data = 24'h2bd4c6;
          13'h0B69 : pic_data = 24'h2bd6d6;
          13'h0B6A : pic_data = 24'h2bc7d4;
          13'h0B6B : pic_data = 24'h2bc0d4;
          13'h0B6C : pic_data = 24'h2bb2d4;
          13'h0B6D : pic_data = 24'h2ba5d4;
          13'h0B6E : pic_data = 24'h2ba2d4;
          13'h0B6F : pic_data = 24'h2b95d4;
          13'h0B70 : pic_data = 24'h2b8dd4;
          13'h0B71 : pic_data = 24'h2b7fd4;
          13'h0B72 : pic_data = 24'h2b73d4;
          13'h0B73 : pic_data = 24'h2b70d4;
          13'h0B74 : pic_data = 24'h2b62d4;
          13'h0B75 : pic_data = 24'h2b5cd4;
          13'h0B76 : pic_data = 24'h2b4cd4;
          13'h0B77 : pic_data = 24'h2b41d4;
          13'h0B78 : pic_data = 24'h2b3cd4;
          13'h0B79 : pic_data = 24'h2b30d4;
          13'h0B7A : pic_data = 24'h2d2ad4;
          13'h0B7B : pic_data = 24'h3c2bd4;
          13'h0B7C : pic_data = 24'h472bd4;
          13'h0B7D : pic_data = 24'h4e2bd4;
          13'h0B7E : pic_data = 24'h5f2bd4;
          13'h0B7F : pic_data = 24'h5e2bd4;
          13'h0B80 : pic_data = 24'h6f2bd4;
          13'h0B81 : pic_data = 24'h7a2bd4;
          13'h0B82 : pic_data = 24'h812bd4;
          13'h0B83 : pic_data = 24'h922bd4;
          13'h0B84 : pic_data = 24'h912bd4;
          13'h0B85 : pic_data = 24'ha22bd4;
          13'h0B86 : pic_data = 24'hab2bd4;
          13'h0B87 : pic_data = 24'hb42bd4;
          13'h0B88 : pic_data = 24'hc52bd4;
          13'h0B89 : pic_data = 24'hc22bd4;
          13'h0B8A : pic_data = 24'hd62bd5;
          13'h0B8B : pic_data = 24'hd42bca;
          13'h0B8C : pic_data = 24'hd42bc3;
          13'h0B8D : pic_data = 24'hd42bb1;
          13'h0B8E : pic_data = 24'hd42ba9;
          13'h0B8F : pic_data = 24'hd42ba1;
          13'h0B90 : pic_data = 24'hd42b98;
          13'h0B91 : pic_data = 24'hd42b90;
          13'h0B92 : pic_data = 24'hd42b7f;
          13'h0B93 : pic_data = 24'hd42b76;
          13'h0B94 : pic_data = 24'hd42b6f;
          13'h0B95 : pic_data = 24'hd42b66;
          13'h0B96 : pic_data = 24'hd42b5f;
          13'h0B97 : pic_data = 24'hd42b4c;
          13'h0B98 : pic_data = 24'hd42b44;
          13'h0B99 : pic_data = 24'hd42b3b;
          13'h0B9A : pic_data = 24'hd5292a;
          13'h0B9B : pic_data = 24'hd5322a;
          13'h0B9C : pic_data = 24'hd53a2a;
          13'h0B9D : pic_data = 24'hd54e2a;
          13'h0B9E : pic_data = 24'hd5542a;
          13'h0B9F : pic_data = 24'hd55e2a;
          13'h0BA0 : pic_data = 24'hd5652a;
          13'h0BA1 : pic_data = 24'hd56e2a;
          13'h0BA2 : pic_data = 24'hd57f2a;
          13'h0BA3 : pic_data = 24'hd5882a;
          13'h0BA4 : pic_data = 24'hd5912a;
          13'h0BA5 : pic_data = 24'hd5982a;
          13'h0BA6 : pic_data = 24'hd5a12a;
          13'h0BA7 : pic_data = 24'hd5b32a;
          13'h0BA8 : pic_data = 24'hd5b92a;
          13'h0BA9 : pic_data = 24'hd5c42a;
          13'h0BAA : pic_data = 24'hd5ca2a;
          13'h0BAB : pic_data = 24'hd7d62a;
          13'h0BAC : pic_data = 24'hc5d52a;
          13'h0BAD : pic_data = 24'hbdd52a;
          13'h0BAE : pic_data = 24'hb3d52a;
          13'h0BAF : pic_data = 24'ha2d52a;
          13'h0BB0 : pic_data = 24'ha3d52a;
          13'h0BB1 : pic_data = 24'h92d52a;
          13'h0BB2 : pic_data = 24'h8bd52a;
          13'h0BB3 : pic_data = 24'h80d52a;
          13'h0BB4 : pic_data = 24'h6fd52a;
          13'h0BB5 : pic_data = 24'h70d52a;
          13'h0BB6 : pic_data = 24'h5fd52a;
          13'h0BB7 : pic_data = 24'h58d52a;
          13'h0BB8 : pic_data = 24'h4dd52a;
          13'h0BB9 : pic_data = 24'h3dd52a;
          13'h0BBA : pic_data = 24'h3dd52a;
          13'h0BBB : pic_data = 24'h2cd52a;
          13'h0BBC : pic_data = 24'h2ad530;
          13'h0BBD : pic_data = 24'h2ad53b;
          13'h0BBE : pic_data = 24'h2ad54a;
          13'h0BBF : pic_data = 24'h2ad551;
          13'h0BC0 : pic_data = 24'h2ad55e;
          13'h0BC1 : pic_data = 24'h2ad562;
          13'h0BC2 : pic_data = 24'h2ad56e;
          13'h0BC3 : pic_data = 24'h2ad57c;
          13'h0BC4 : pic_data = 24'h2ad584;
          13'h0BC5 : pic_data = 24'h2ad591;
          13'h0BC6 : pic_data = 24'h2ad595;
          13'h0BC7 : pic_data = 24'h2ad5a1;
          13'h0BC8 : pic_data = 24'h2ad5af;
          13'h0BC9 : pic_data = 24'h2ad5b6;
          13'h0BCA : pic_data = 24'h2ad5c5;
          13'h0BCB : pic_data = 24'h2ad5c7;
          13'h0BCC : pic_data = 24'h2ad6d6;
          13'h0BCD : pic_data = 24'h2ac7d5;
          13'h0BCE : pic_data = 24'h2ac0d5;
          13'h0BCF : pic_data = 24'h2ab2d5;
          13'h0BD0 : pic_data = 24'h2aa6d5;
          13'h0BD1 : pic_data = 24'h2aa2d5;
          13'h0BD2 : pic_data = 24'h2a95d5;
          13'h0BD3 : pic_data = 24'h2a8dd5;
          13'h0BD4 : pic_data = 24'h2a7fd5;
          13'h0BD5 : pic_data = 24'h2a73d5;
          13'h0BD6 : pic_data = 24'h2a6fd5;
          13'h0BD7 : pic_data = 24'h2a62d5;
          13'h0BD8 : pic_data = 24'h2a5bd5;
          13'h0BD9 : pic_data = 24'h2a4cd5;
          13'h0BDA : pic_data = 24'h2a41d5;
          13'h0BDB : pic_data = 24'h2a3cd5;
          13'h0BDC : pic_data = 24'h2a30d5;
          13'h0BDD : pic_data = 24'h2c2ad5;
          13'h0BDE : pic_data = 24'h3c2ad5;
          13'h0BDF : pic_data = 24'h472ad5;
          13'h0BE0 : pic_data = 24'h4e2ad5;
          13'h0BE1 : pic_data = 24'h5f2ad5;
          13'h0BE2 : pic_data = 24'h5e2ad5;
          13'h0BE3 : pic_data = 24'h6f2ad5;
          13'h0BE4 : pic_data = 24'h7a2ad5;
          13'h0BE5 : pic_data = 24'h812ad5;
          13'h0BE6 : pic_data = 24'h922ad5;
          13'h0BE7 : pic_data = 24'h912ad5;
          13'h0BE8 : pic_data = 24'ha22ad5;
          13'h0BE9 : pic_data = 24'hac2ad5;
          13'h0BEA : pic_data = 24'hb42ad5;
          13'h0BEB : pic_data = 24'hc52ad5;
          13'h0BEC : pic_data = 24'hc32ad5;
          13'h0BED : pic_data = 24'hd72ad6;
          13'h0BEE : pic_data = 24'hd52aca;
          13'h0BEF : pic_data = 24'hd52ac4;
          13'h0BF0 : pic_data = 24'hd52ab2;
          13'h0BF1 : pic_data = 24'hd52aa9;
          13'h0BF2 : pic_data = 24'hd52aa2;
          13'h0BF3 : pic_data = 24'hd52a99;
          13'h0BF4 : pic_data = 24'hd52a90;
          13'h0BF5 : pic_data = 24'hd52a7f;
          13'h0BF6 : pic_data = 24'hd52a76;
          13'h0BF7 : pic_data = 24'hd52a6f;
          13'h0BF8 : pic_data = 24'hd52a65;
          13'h0BF9 : pic_data = 24'hd52a5f;
          13'h0BFA : pic_data = 24'hd52a4b;
          13'h0BFB : pic_data = 24'hd52a43;
          13'h0BFC : pic_data = 24'hd52a3a;
          13'h0BFD : pic_data = 24'hd32b2c;
          13'h0BFE : pic_data = 24'hd3332c;
          13'h0BFF : pic_data = 24'hd33b2c;
          13'h0C00 : pic_data = 24'hd34e2c;
          13'h0C01 : pic_data = 24'hd3552c;
          13'h0C02 : pic_data = 24'hd35e2c;
          13'h0C03 : pic_data = 24'hd3662c;
          13'h0C04 : pic_data = 24'hd36e2c;
          13'h0C05 : pic_data = 24'hd37f2c;
          13'h0C06 : pic_data = 24'hd3872c;
          13'h0C07 : pic_data = 24'hd3902c;
          13'h0C08 : pic_data = 24'hd3982c;
          13'h0C09 : pic_data = 24'hd3a02c;
          13'h0C0A : pic_data = 24'hd3b22c;
          13'h0C0B : pic_data = 24'hd3b92c;
          13'h0C0C : pic_data = 24'hd3c32c;
          13'h0C0D : pic_data = 24'hd3c92c;
          13'h0C0E : pic_data = 24'hd5d42c;
          13'h0C0F : pic_data = 24'hc3d32c;
          13'h0C10 : pic_data = 24'hbcd32c;
          13'h0C11 : pic_data = 24'hb2d32c;
          13'h0C12 : pic_data = 24'ha1d32c;
          13'h0C13 : pic_data = 24'ha2d32c;
          13'h0C14 : pic_data = 24'h91d32c;
          13'h0C15 : pic_data = 24'h8ad32c;
          13'h0C16 : pic_data = 24'h80d32c;
          13'h0C17 : pic_data = 24'h6fd32c;
          13'h0C18 : pic_data = 24'h70d32c;
          13'h0C19 : pic_data = 24'h5fd32c;
          13'h0C1A : pic_data = 24'h58d32c;
          13'h0C1B : pic_data = 24'h4dd32c;
          13'h0C1C : pic_data = 24'h3ed32c;
          13'h0C1D : pic_data = 24'h3ed32c;
          13'h0C1E : pic_data = 24'h2dd32b;
          13'h0C1F : pic_data = 24'h2bd331;
          13'h0C20 : pic_data = 24'h2cd33c;
          13'h0C21 : pic_data = 24'h2cd34b;
          13'h0C22 : pic_data = 24'h2cd352;
          13'h0C23 : pic_data = 24'h2cd35f;
          13'h0C24 : pic_data = 24'h2cd362;
          13'h0C25 : pic_data = 24'h2cd36f;
          13'h0C26 : pic_data = 24'h2cd37c;
          13'h0C27 : pic_data = 24'h2cd384;
          13'h0C28 : pic_data = 24'h2cd391;
          13'h0C29 : pic_data = 24'h2cd394;
          13'h0C2A : pic_data = 24'h2cd3a1;
          13'h0C2B : pic_data = 24'h2cd3ae;
          13'h0C2C : pic_data = 24'h2cd3b5;
          13'h0C2D : pic_data = 24'h2cd3c4;
          13'h0C2E : pic_data = 24'h2cd3c5;
          13'h0C2F : pic_data = 24'h2cd5d5;
          13'h0C30 : pic_data = 24'h2cc6d3;
          13'h0C31 : pic_data = 24'h2cbfd3;
          13'h0C32 : pic_data = 24'h2cb2d3;
          13'h0C33 : pic_data = 24'h2ca5d3;
          13'h0C34 : pic_data = 24'h2ca2d3;
          13'h0C35 : pic_data = 24'h2c95d3;
          13'h0C36 : pic_data = 24'h2c8dd3;
          13'h0C37 : pic_data = 24'h2c7fd3;
          13'h0C38 : pic_data = 24'h2c73d3;
          13'h0C39 : pic_data = 24'h2c70d3;
          13'h0C3A : pic_data = 24'h2c63d3;
          13'h0C3B : pic_data = 24'h2c5cd3;
          13'h0C3C : pic_data = 24'h2c4dd3;
          13'h0C3D : pic_data = 24'h2c41d3;
          13'h0C3E : pic_data = 24'h2c3dd3;
          13'h0C3F : pic_data = 24'h2b31d3;
          13'h0C40 : pic_data = 24'h2d2bd3;
          13'h0C41 : pic_data = 24'h3d2cd3;
          13'h0C42 : pic_data = 24'h472cd3;
          13'h0C43 : pic_data = 24'h4e2cd3;
          13'h0C44 : pic_data = 24'h602cd3;
          13'h0C45 : pic_data = 24'h5e2cd3;
          13'h0C46 : pic_data = 24'h6f2cd3;
          13'h0C47 : pic_data = 24'h7a2cd3;
          13'h0C48 : pic_data = 24'h812cd3;
          13'h0C49 : pic_data = 24'h922cd3;
          13'h0C4A : pic_data = 24'h902cd3;
          13'h0C4B : pic_data = 24'ha12cd3;
          13'h0C4C : pic_data = 24'hab2cd3;
          13'h0C4D : pic_data = 24'hb32cd3;
          13'h0C4E : pic_data = 24'hc42cd3;
          13'h0C4F : pic_data = 24'hc22cd3;
          13'h0C50 : pic_data = 24'hd52cd4;
          13'h0C51 : pic_data = 24'hd32cc9;
          13'h0C52 : pic_data = 24'hd32cc2;
          13'h0C53 : pic_data = 24'hd32cb1;
          13'h0C54 : pic_data = 24'hd32ca9;
          13'h0C55 : pic_data = 24'hd32ca1;
          13'h0C56 : pic_data = 24'hd32c98;
          13'h0C57 : pic_data = 24'hd32c90;
          13'h0C58 : pic_data = 24'hd32c7f;
          13'h0C59 : pic_data = 24'hd32c76;
          13'h0C5A : pic_data = 24'hd32c6f;
          13'h0C5B : pic_data = 24'hd32c66;
          13'h0C5C : pic_data = 24'hd32c5f;
          13'h0C5D : pic_data = 24'hd32c4c;
          13'h0C5E : pic_data = 24'hd32c44;
          13'h0C5F : pic_data = 24'hd32c3b;
          13'h0C60 : pic_data = 24'hcf2e2f;
          13'h0C61 : pic_data = 24'hcf372f;
          13'h0C62 : pic_data = 24'hcf3e2f;
          13'h0C63 : pic_data = 24'hcf502f;
          13'h0C64 : pic_data = 24'hcf572f;
          13'h0C65 : pic_data = 24'hcf602f;
          13'h0C66 : pic_data = 24'hcf662f;
          13'h0C67 : pic_data = 24'hcf6f2f;
          13'h0C68 : pic_data = 24'hcf7f2f;
          13'h0C69 : pic_data = 24'hcf862f;
          13'h0C6A : pic_data = 24'hcf8e2f;
          13'h0C6B : pic_data = 24'hcf952f;
          13'h0C6C : pic_data = 24'hcf9d2f;
          13'h0C6D : pic_data = 24'hcfaf2f;
          13'h0C6E : pic_data = 24'hcfb62f;
          13'h0C6F : pic_data = 24'hcfbf2f;
          13'h0C70 : pic_data = 24'hcfc62f;
          13'h0C71 : pic_data = 24'hd1d02f;
          13'h0C72 : pic_data = 24'hbfcf2f;
          13'h0C73 : pic_data = 24'hbacf2f;
          13'h0C74 : pic_data = 24'hb0cf2f;
          13'h0C75 : pic_data = 24'h9fcf2f;
          13'h0C76 : pic_data = 24'ha0cf2f;
          13'h0C77 : pic_data = 24'h90cf2f;
          13'h0C78 : pic_data = 24'h88cf2f;
          13'h0C79 : pic_data = 24'h80cf2f;
          13'h0C7A : pic_data = 24'h70cf2f;
          13'h0C7B : pic_data = 24'h71cf2f;
          13'h0C7C : pic_data = 24'h61cf2f;
          13'h0C7D : pic_data = 24'h5acf2f;
          13'h0C7E : pic_data = 24'h4fcf2f;
          13'h0C7F : pic_data = 24'h41cf2f;
          13'h0C80 : pic_data = 24'h40cf2f;
          13'h0C81 : pic_data = 24'h31cf2e;
          13'h0C82 : pic_data = 24'h2ecf33;
          13'h0C83 : pic_data = 24'h2fcf3f;
          13'h0C84 : pic_data = 24'h2fcf4c;
          13'h0C85 : pic_data = 24'h2fcf53;
          13'h0C86 : pic_data = 24'h2fcf61;
          13'h0C87 : pic_data = 24'h2fcf64;
          13'h0C88 : pic_data = 24'h2fcf6f;
          13'h0C89 : pic_data = 24'h2fcf7d;
          13'h0C8A : pic_data = 24'h2fcf83;
          13'h0C8B : pic_data = 24'h2fcf8f;
          13'h0C8C : pic_data = 24'h2fcf91;
          13'h0C8D : pic_data = 24'h2fcf9e;
          13'h0C8E : pic_data = 24'h2fcfac;
          13'h0C8F : pic_data = 24'h2fcfb3;
          13'h0C90 : pic_data = 24'h2fcfc0;
          13'h0C91 : pic_data = 24'h2fcfc2;
          13'h0C92 : pic_data = 24'h2fd1d1;
          13'h0C93 : pic_data = 24'h2fc3cf;
          13'h0C94 : pic_data = 24'h2fbccf;
          13'h0C95 : pic_data = 24'h2fafcf;
          13'h0C96 : pic_data = 24'h2fa2cf;
          13'h0C97 : pic_data = 24'h2f9fcf;
          13'h0C98 : pic_data = 24'h2f93cf;
          13'h0C99 : pic_data = 24'h2f8ccf;
          13'h0C9A : pic_data = 24'h2f7fcf;
          13'h0C9B : pic_data = 24'h2f74cf;
          13'h0C9C : pic_data = 24'h2f70cf;
          13'h0C9D : pic_data = 24'h2f64cf;
          13'h0C9E : pic_data = 24'h2f5dcf;
          13'h0C9F : pic_data = 24'h2f4ecf;
          13'h0CA0 : pic_data = 24'h2f43cf;
          13'h0CA1 : pic_data = 24'h2f40cf;
          13'h0CA2 : pic_data = 24'h2e33cf;
          13'h0CA3 : pic_data = 24'h312ecf;
          13'h0CA4 : pic_data = 24'h3f2fcf;
          13'h0CA5 : pic_data = 24'h492fcf;
          13'h0CA6 : pic_data = 24'h502fcf;
          13'h0CA7 : pic_data = 24'h612fcf;
          13'h0CA8 : pic_data = 24'h602fcf;
          13'h0CA9 : pic_data = 24'h702fcf;
          13'h0CAA : pic_data = 24'h7a2fcf;
          13'h0CAB : pic_data = 24'h812fcf;
          13'h0CAC : pic_data = 24'h902fcf;
          13'h0CAD : pic_data = 24'h8f2fcf;
          13'h0CAE : pic_data = 24'h9f2fcf;
          13'h0CAF : pic_data = 24'ha82fcf;
          13'h0CB0 : pic_data = 24'haf2fcf;
          13'h0CB1 : pic_data = 24'hc12fcf;
          13'h0CB2 : pic_data = 24'hbe2fcf;
          13'h0CB3 : pic_data = 24'hd12fd0;
          13'h0CB4 : pic_data = 24'hcf2fc6;
          13'h0CB5 : pic_data = 24'hcf2fbf;
          13'h0CB6 : pic_data = 24'hcf2fae;
          13'h0CB7 : pic_data = 24'hcf2fa6;
          13'h0CB8 : pic_data = 24'hcf2f9e;
          13'h0CB9 : pic_data = 24'hcf2f95;
          13'h0CBA : pic_data = 24'hcf2f8e;
          13'h0CBB : pic_data = 24'hcf2f7f;
          13'h0CBC : pic_data = 24'hcf2f76;
          13'h0CBD : pic_data = 24'hcf2f70;
          13'h0CBE : pic_data = 24'hcf2f68;
          13'h0CBF : pic_data = 24'hcf2f61;
          13'h0CC0 : pic_data = 24'hcf2f4e;
          13'h0CC1 : pic_data = 24'hcf2f47;
          13'h0CC2 : pic_data = 24'hcf2f3e;
          13'h0CC3 : pic_data = 24'hd02d2e;
          13'h0CC4 : pic_data = 24'hd0362e;
          13'h0CC5 : pic_data = 24'hd03d2e;
          13'h0CC6 : pic_data = 24'hd04f2e;
          13'h0CC7 : pic_data = 24'hd0562e;
          13'h0CC8 : pic_data = 24'hd0602e;
          13'h0CC9 : pic_data = 24'hd0662e;
          13'h0CCA : pic_data = 24'hd06f2e;
          13'h0CCB : pic_data = 24'hd07f2e;
          13'h0CCC : pic_data = 24'hd0872e;
          13'h0CCD : pic_data = 24'hd08f2e;
          13'h0CCE : pic_data = 24'hd0952e;
          13'h0CCF : pic_data = 24'hd09e2e;
          13'h0CD0 : pic_data = 24'hd0b02e;
          13'h0CD1 : pic_data = 24'hd0b72e;
          13'h0CD2 : pic_data = 24'hd0c02e;
          13'h0CD3 : pic_data = 24'hd0c72e;
          13'h0CD4 : pic_data = 24'hd2d12e;
          13'h0CD5 : pic_data = 24'hc0d02e;
          13'h0CD6 : pic_data = 24'hbad02e;
          13'h0CD7 : pic_data = 24'hb0d02e;
          13'h0CD8 : pic_data = 24'h9fd02e;
          13'h0CD9 : pic_data = 24'ha0d02e;
          13'h0CDA : pic_data = 24'h90d02e;
          13'h0CDB : pic_data = 24'h89d02e;
          13'h0CDC : pic_data = 24'h80d02e;
          13'h0CDD : pic_data = 24'h70d02e;
          13'h0CDE : pic_data = 24'h71d02e;
          13'h0CDF : pic_data = 24'h61d02e;
          13'h0CE0 : pic_data = 24'h5ad02e;
          13'h0CE1 : pic_data = 24'h4ed02e;
          13'h0CE2 : pic_data = 24'h40d02e;
          13'h0CE3 : pic_data = 24'h3fd02e;
          13'h0CE4 : pic_data = 24'h30d02d;
          13'h0CE5 : pic_data = 24'h2ed032;
          13'h0CE6 : pic_data = 24'h2ed03e;
          13'h0CE7 : pic_data = 24'h2ed04c;
          13'h0CE8 : pic_data = 24'h2ed053;
          13'h0CE9 : pic_data = 24'h2ed060;
          13'h0CEA : pic_data = 24'h2ed064;
          13'h0CEB : pic_data = 24'h2ed06f;
          13'h0CEC : pic_data = 24'h2ed07d;
          13'h0CED : pic_data = 24'h2ed083;
          13'h0CEE : pic_data = 24'h2ed08f;
          13'h0CEF : pic_data = 24'h2ed092;
          13'h0CF0 : pic_data = 24'h2ed09e;
          13'h0CF1 : pic_data = 24'h2ed0ac;
          13'h0CF2 : pic_data = 24'h2ed0b3;
          13'h0CF3 : pic_data = 24'h2ed0c1;
          13'h0CF4 : pic_data = 24'h2ed0c3;
          13'h0CF5 : pic_data = 24'h2ed1d1;
          13'h0CF6 : pic_data = 24'h2ec3d0;
          13'h0CF7 : pic_data = 24'h2ebcd0;
          13'h0CF8 : pic_data = 24'h2eb0d0;
          13'h0CF9 : pic_data = 24'h2ea3d0;
          13'h0CFA : pic_data = 24'h2e9fd0;
          13'h0CFB : pic_data = 24'h2e93d0;
          13'h0CFC : pic_data = 24'h2e8cd0;
          13'h0CFD : pic_data = 24'h2e7fd0;
          13'h0CFE : pic_data = 24'h2e74d0;
          13'h0CFF : pic_data = 24'h2e70d0;
          13'h0D00 : pic_data = 24'h2e64d0;
          13'h0D01 : pic_data = 24'h2e5dd0;
          13'h0D02 : pic_data = 24'h2e4ed0;
          13'h0D03 : pic_data = 24'h2e42d0;
          13'h0D04 : pic_data = 24'h2e3fd0;
          13'h0D05 : pic_data = 24'h2e32d0;
          13'h0D06 : pic_data = 24'h302dd0;
          13'h0D07 : pic_data = 24'h3f2ed0;
          13'h0D08 : pic_data = 24'h482ed0;
          13'h0D09 : pic_data = 24'h4f2ed0;
          13'h0D0A : pic_data = 24'h612ed0;
          13'h0D0B : pic_data = 24'h602ed0;
          13'h0D0C : pic_data = 24'h702ed0;
          13'h0D0D : pic_data = 24'h7a2ed0;
          13'h0D0E : pic_data = 24'h812ed0;
          13'h0D0F : pic_data = 24'h902ed0;
          13'h0D10 : pic_data = 24'h8f2ed0;
          13'h0D11 : pic_data = 24'h9f2ed0;
          13'h0D12 : pic_data = 24'ha92ed0;
          13'h0D13 : pic_data = 24'hb02ed0;
          13'h0D14 : pic_data = 24'hc22ed0;
          13'h0D15 : pic_data = 24'hbf2ed0;
          13'h0D16 : pic_data = 24'hd22ed1;
          13'h0D17 : pic_data = 24'hd02ec7;
          13'h0D18 : pic_data = 24'hd02ec0;
          13'h0D19 : pic_data = 24'hd02eaf;
          13'h0D1A : pic_data = 24'hd02ea7;
          13'h0D1B : pic_data = 24'hd02e9f;
          13'h0D1C : pic_data = 24'hd02e95;
          13'h0D1D : pic_data = 24'hd02e8e;
          13'h0D1E : pic_data = 24'hd02e7f;
          13'h0D1F : pic_data = 24'hd02e76;
          13'h0D20 : pic_data = 24'hd02e70;
          13'h0D21 : pic_data = 24'hd02e67;
          13'h0D22 : pic_data = 24'hd02e61;
          13'h0D23 : pic_data = 24'hd02e4d;
          13'h0D24 : pic_data = 24'hd02e46;
          13'h0D25 : pic_data = 24'hd02e3d;
          13'h0D26 : pic_data = 24'hcc3132;
          13'h0D27 : pic_data = 24'hcc3932;
          13'h0D28 : pic_data = 24'hcc4032;
          13'h0D29 : pic_data = 24'hcc5232;
          13'h0D2A : pic_data = 24'hcc5832;
          13'h0D2B : pic_data = 24'hcc6132;
          13'h0D2C : pic_data = 24'hcc6732;
          13'h0D2D : pic_data = 24'hcc7032;
          13'h0D2E : pic_data = 24'hcc7f32;
          13'h0D2F : pic_data = 24'hcc8632;
          13'h0D30 : pic_data = 24'hcc8e32;
          13'h0D31 : pic_data = 24'hcc9432;
          13'h0D32 : pic_data = 24'hcc9d32;
          13'h0D33 : pic_data = 24'hccad32;
          13'h0D34 : pic_data = 24'hccb432;
          13'h0D35 : pic_data = 24'hccbd32;
          13'h0D36 : pic_data = 24'hccc332;
          13'h0D37 : pic_data = 24'hcecd32;
          13'h0D38 : pic_data = 24'hbdcc32;
          13'h0D39 : pic_data = 24'hb7cc32;
          13'h0D3A : pic_data = 24'hadcc32;
          13'h0D3B : pic_data = 24'h9ecc32;
          13'h0D3C : pic_data = 24'h9fcc32;
          13'h0D3D : pic_data = 24'h8fcc32;
          13'h0D3E : pic_data = 24'h89cc32;
          13'h0D3F : pic_data = 24'h80cc32;
          13'h0D40 : pic_data = 24'h71cc32;
          13'h0D41 : pic_data = 24'h72cc32;
          13'h0D42 : pic_data = 24'h62cc32;
          13'h0D43 : pic_data = 24'h5ccc32;
          13'h0D44 : pic_data = 24'h51cc32;
          13'h0D45 : pic_data = 24'h43cc32;
          13'h0D46 : pic_data = 24'h42cc32;
          13'h0D47 : pic_data = 24'h34cc31;
          13'h0D48 : pic_data = 24'h32cc36;
          13'h0D49 : pic_data = 24'h32cc41;
          13'h0D4A : pic_data = 24'h32cc4f;
          13'h0D4B : pic_data = 24'h32cc56;
          13'h0D4C : pic_data = 24'h32cc61;
          13'h0D4D : pic_data = 24'h32cc65;
          13'h0D4E : pic_data = 24'h32cc70;
          13'h0D4F : pic_data = 24'h32cc7d;
          13'h0D50 : pic_data = 24'h32cc83;
          13'h0D51 : pic_data = 24'h32cc8e;
          13'h0D52 : pic_data = 24'h32cc91;
          13'h0D53 : pic_data = 24'h32cc9e;
          13'h0D54 : pic_data = 24'h32cca9;
          13'h0D55 : pic_data = 24'h32ccb0;
          13'h0D56 : pic_data = 24'h32ccbe;
          13'h0D57 : pic_data = 24'h32ccc0;
          13'h0D58 : pic_data = 24'h32cdcd;
          13'h0D59 : pic_data = 24'h32c1cc;
          13'h0D5A : pic_data = 24'h32b9cc;
          13'h0D5B : pic_data = 24'h32adcc;
          13'h0D5C : pic_data = 24'h32a1cc;
          13'h0D5D : pic_data = 24'h329ecc;
          13'h0D5E : pic_data = 24'h3292cc;
          13'h0D5F : pic_data = 24'h328bcc;
          13'h0D60 : pic_data = 24'h327fcc;
          13'h0D61 : pic_data = 24'h3274cc;
          13'h0D62 : pic_data = 24'h3271cc;
          13'h0D63 : pic_data = 24'h3265cc;
          13'h0D64 : pic_data = 24'h325ecc;
          13'h0D65 : pic_data = 24'h3251cc;
          13'h0D66 : pic_data = 24'h3245cc;
          13'h0D67 : pic_data = 24'h3242cc;
          13'h0D68 : pic_data = 24'h3236cc;
          13'h0D69 : pic_data = 24'h3331cc;
          13'h0D6A : pic_data = 24'h4132cc;
          13'h0D6B : pic_data = 24'h4b32cc;
          13'h0D6C : pic_data = 24'h5232cc;
          13'h0D6D : pic_data = 24'h6232cc;
          13'h0D6E : pic_data = 24'h6132cc;
          13'h0D6F : pic_data = 24'h7132cc;
          13'h0D70 : pic_data = 24'h7a32cc;
          13'h0D71 : pic_data = 24'h8132cc;
          13'h0D72 : pic_data = 24'h8f32cc;
          13'h0D73 : pic_data = 24'h8e32cc;
          13'h0D74 : pic_data = 24'h9e32cc;
          13'h0D75 : pic_data = 24'ha732cc;
          13'h0D76 : pic_data = 24'had32cc;
          13'h0D77 : pic_data = 24'hbf32cc;
          13'h0D78 : pic_data = 24'hbc32cc;
          13'h0D79 : pic_data = 24'hce32cd;
          13'h0D7A : pic_data = 24'hcc32c3;
          13'h0D7B : pic_data = 24'hcc32bd;
          13'h0D7C : pic_data = 24'hcc32ac;
          13'h0D7D : pic_data = 24'hcc32a5;
          13'h0D7E : pic_data = 24'hcc329e;
          13'h0D7F : pic_data = 24'hcc3295;
          13'h0D80 : pic_data = 24'hcc328d;
          13'h0D81 : pic_data = 24'hcc327f;
          13'h0D82 : pic_data = 24'hcc3277;
          13'h0D83 : pic_data = 24'hcc3270;
          13'h0D84 : pic_data = 24'hcc3268;
          13'h0D85 : pic_data = 24'hcc3261;
          13'h0D86 : pic_data = 24'hcc3250;
          13'h0D87 : pic_data = 24'hcc3249;
          13'h0D88 : pic_data = 24'hcc3240;
          13'h0D89 : pic_data = 24'hcb3233;
          13'h0D8A : pic_data = 24'hcb3933;
          13'h0D8B : pic_data = 24'hcb4133;
          13'h0D8C : pic_data = 24'hcb5333;
          13'h0D8D : pic_data = 24'hcb5833;
          13'h0D8E : pic_data = 24'hcb6133;
          13'h0D8F : pic_data = 24'hcb6733;
          13'h0D90 : pic_data = 24'hcb7033;
          13'h0D91 : pic_data = 24'hcb7f33;
          13'h0D92 : pic_data = 24'hcb8533;
          13'h0D93 : pic_data = 24'hcb8e33;
          13'h0D94 : pic_data = 24'hcb9433;
          13'h0D95 : pic_data = 24'hcb9d33;
          13'h0D96 : pic_data = 24'hcbac33;
          13'h0D97 : pic_data = 24'hcbb333;
          13'h0D98 : pic_data = 24'hcbbd33;
          13'h0D99 : pic_data = 24'hcbc233;
          13'h0D9A : pic_data = 24'hcdcd33;
          13'h0D9B : pic_data = 24'hbdcb33;
          13'h0D9C : pic_data = 24'hb7cb33;
          13'h0D9D : pic_data = 24'hadcb33;
          13'h0D9E : pic_data = 24'h9ecb33;
          13'h0D9F : pic_data = 24'h9fcb33;
          13'h0DA0 : pic_data = 24'h8fcb33;
          13'h0DA1 : pic_data = 24'h89cb33;
          13'h0DA2 : pic_data = 24'h80cb33;
          13'h0DA3 : pic_data = 24'h71cb33;
          13'h0DA4 : pic_data = 24'h72cb33;
          13'h0DA5 : pic_data = 24'h62cb33;
          13'h0DA6 : pic_data = 24'h5ccb33;
          13'h0DA7 : pic_data = 24'h52cb33;
          13'h0DA8 : pic_data = 24'h43cb33;
          13'h0DA9 : pic_data = 24'h43cb33;
          13'h0DAA : pic_data = 24'h34cb32;
          13'h0DAB : pic_data = 24'h32cb37;
          13'h0DAC : pic_data = 24'h33cb41;
          13'h0DAD : pic_data = 24'h33cb4f;
          13'h0DAE : pic_data = 24'h33cb56;
          13'h0DAF : pic_data = 24'h33cb61;
          13'h0DB0 : pic_data = 24'h33cb65;
          13'h0DB1 : pic_data = 24'h33cb70;
          13'h0DB2 : pic_data = 24'h33cb7d;
          13'h0DB3 : pic_data = 24'h33cb83;
          13'h0DB4 : pic_data = 24'h33cb8e;
          13'h0DB5 : pic_data = 24'h33cb90;
          13'h0DB6 : pic_data = 24'h33cb9e;
          13'h0DB7 : pic_data = 24'h33cba9;
          13'h0DB8 : pic_data = 24'h33cbb0;
          13'h0DB9 : pic_data = 24'h33cbbd;
          13'h0DBA : pic_data = 24'h33cbc0;
          13'h0DBB : pic_data = 24'h33cdcd;
          13'h0DBC : pic_data = 24'h33c0cb;
          13'h0DBD : pic_data = 24'h33b9cb;
          13'h0DBE : pic_data = 24'h33accb;
          13'h0DBF : pic_data = 24'h33a1cb;
          13'h0DC0 : pic_data = 24'h339ecb;
          13'h0DC1 : pic_data = 24'h3392cb;
          13'h0DC2 : pic_data = 24'h338bcb;
          13'h0DC3 : pic_data = 24'h3380cb;
          13'h0DC4 : pic_data = 24'h3374cb;
          13'h0DC5 : pic_data = 24'h3371cb;
          13'h0DC6 : pic_data = 24'h3365cb;
          13'h0DC7 : pic_data = 24'h335ecb;
          13'h0DC8 : pic_data = 24'h3351cb;
          13'h0DC9 : pic_data = 24'h3346cb;
          13'h0DCA : pic_data = 24'h3342cb;
          13'h0DCB : pic_data = 24'h3237cb;
          13'h0DCC : pic_data = 24'h3332cb;
          13'h0DCD : pic_data = 24'h4233cb;
          13'h0DCE : pic_data = 24'h4c33cb;
          13'h0DCF : pic_data = 24'h5333cb;
          13'h0DD0 : pic_data = 24'h6233cb;
          13'h0DD1 : pic_data = 24'h6133cb;
          13'h0DD2 : pic_data = 24'h7133cb;
          13'h0DD3 : pic_data = 24'h7a33cb;
          13'h0DD4 : pic_data = 24'h8133cb;
          13'h0DD5 : pic_data = 24'h8f33cb;
          13'h0DD6 : pic_data = 24'h8e33cb;
          13'h0DD7 : pic_data = 24'h9e33cb;
          13'h0DD8 : pic_data = 24'ha733cb;
          13'h0DD9 : pic_data = 24'hac33cb;
          13'h0DDA : pic_data = 24'hbe33cb;
          13'h0DDB : pic_data = 24'hbc33cb;
          13'h0DDC : pic_data = 24'hcd33cd;
          13'h0DDD : pic_data = 24'hcb33c2;
          13'h0DDE : pic_data = 24'hcb33bc;
          13'h0DDF : pic_data = 24'hcb33ac;
          13'h0DE0 : pic_data = 24'hcb33a4;
          13'h0DE1 : pic_data = 24'hcb339e;
          13'h0DE2 : pic_data = 24'hcb3394;
          13'h0DE3 : pic_data = 24'hcb338d;
          13'h0DE4 : pic_data = 24'hcb337f;
          13'h0DE5 : pic_data = 24'hcb3377;
          13'h0DE6 : pic_data = 24'hcb3371;
          13'h0DE7 : pic_data = 24'hcb3369;
          13'h0DE8 : pic_data = 24'hcb3361;
          13'h0DE9 : pic_data = 24'hcb3351;
          13'h0DEA : pic_data = 24'hcb334a;
          13'h0DEB : pic_data = 24'hcb3341;
          13'h0DEC : pic_data = 24'hcc3132;
          13'h0DED : pic_data = 24'hcc3932;
          13'h0DEE : pic_data = 24'hcc4032;
          13'h0DEF : pic_data = 24'hcc5232;
          13'h0DF0 : pic_data = 24'hcc5832;
          13'h0DF1 : pic_data = 24'hcc6032;
          13'h0DF2 : pic_data = 24'hcc6732;
          13'h0DF3 : pic_data = 24'hcc7032;
          13'h0DF4 : pic_data = 24'hcc7f32;
          13'h0DF5 : pic_data = 24'hcc8532;
          13'h0DF6 : pic_data = 24'hcc8e32;
          13'h0DF7 : pic_data = 24'hcc9432;
          13'h0DF8 : pic_data = 24'hcc9d32;
          13'h0DF9 : pic_data = 24'hccac32;
          13'h0DFA : pic_data = 24'hccb432;
          13'h0DFB : pic_data = 24'hccbd32;
          13'h0DFC : pic_data = 24'hccc332;
          13'h0DFD : pic_data = 24'hcecd32;
          13'h0DFE : pic_data = 24'hbdcc32;
          13'h0DFF : pic_data = 24'hb7cc32;
          13'h0E00 : pic_data = 24'hadcc32;
          13'h0E01 : pic_data = 24'h9ecc32;
          13'h0E02 : pic_data = 24'h9fcc32;
          13'h0E03 : pic_data = 24'h8fcc32;
          13'h0E04 : pic_data = 24'h89cc32;
          13'h0E05 : pic_data = 24'h80cc32;
          13'h0E06 : pic_data = 24'h71cc32;
          13'h0E07 : pic_data = 24'h72cc32;
          13'h0E08 : pic_data = 24'h61cc32;
          13'h0E09 : pic_data = 24'h5ccc32;
          13'h0E0A : pic_data = 24'h52cc32;
          13'h0E0B : pic_data = 24'h43cc32;
          13'h0E0C : pic_data = 24'h42cc32;
          13'h0E0D : pic_data = 24'h34cc31;
          13'h0E0E : pic_data = 24'h32cc36;
          13'h0E0F : pic_data = 24'h32cc41;
          13'h0E10 : pic_data = 24'h32cc4f;
          13'h0E11 : pic_data = 24'h32cc56;
          13'h0E12 : pic_data = 24'h32cc61;
          13'h0E13 : pic_data = 24'h32cc65;
          13'h0E14 : pic_data = 24'h32cc70;
          13'h0E15 : pic_data = 24'h32cc7d;
          13'h0E16 : pic_data = 24'h32cc83;
          13'h0E17 : pic_data = 24'h32cc8e;
          13'h0E18 : pic_data = 24'h32cc91;
          13'h0E19 : pic_data = 24'h32cc9e;
          13'h0E1A : pic_data = 24'h32cca9;
          13'h0E1B : pic_data = 24'h32ccb0;
          13'h0E1C : pic_data = 24'h32ccbe;
          13'h0E1D : pic_data = 24'h32ccc0;
          13'h0E1E : pic_data = 24'h32cdcd;
          13'h0E1F : pic_data = 24'h32c1cc;
          13'h0E20 : pic_data = 24'h32b9cc;
          13'h0E21 : pic_data = 24'h32adcc;
          13'h0E22 : pic_data = 24'h32a1cc;
          13'h0E23 : pic_data = 24'h329fcc;
          13'h0E24 : pic_data = 24'h3292cc;
          13'h0E25 : pic_data = 24'h328bcc;
          13'h0E26 : pic_data = 24'h3280cc;
          13'h0E27 : pic_data = 24'h3274cc;
          13'h0E28 : pic_data = 24'h3271cc;
          13'h0E29 : pic_data = 24'h3265cc;
          13'h0E2A : pic_data = 24'h325ecc;
          13'h0E2B : pic_data = 24'h3251cc;
          13'h0E2C : pic_data = 24'h3245cc;
          13'h0E2D : pic_data = 24'h3242cc;
          13'h0E2E : pic_data = 24'h3236cc;
          13'h0E2F : pic_data = 24'h3331cc;
          13'h0E30 : pic_data = 24'h4132cc;
          13'h0E31 : pic_data = 24'h4b32cc;
          13'h0E32 : pic_data = 24'h5332cc;
          13'h0E33 : pic_data = 24'h6232cc;
          13'h0E34 : pic_data = 24'h6132cc;
          13'h0E35 : pic_data = 24'h7132cc;
          13'h0E36 : pic_data = 24'h7a32cc;
          13'h0E37 : pic_data = 24'h8132cc;
          13'h0E38 : pic_data = 24'h8f32cc;
          13'h0E39 : pic_data = 24'h8e32cc;
          13'h0E3A : pic_data = 24'h9e32cc;
          13'h0E3B : pic_data = 24'ha732cc;
          13'h0E3C : pic_data = 24'had32cc;
          13'h0E3D : pic_data = 24'hbf32cc;
          13'h0E3E : pic_data = 24'hbc32cc;
          13'h0E3F : pic_data = 24'hce32cd;
          13'h0E40 : pic_data = 24'hcc32c3;
          13'h0E41 : pic_data = 24'hcc32bd;
          13'h0E42 : pic_data = 24'hcc32ac;
          13'h0E43 : pic_data = 24'hcc32a5;
          13'h0E44 : pic_data = 24'hcc329e;
          13'h0E45 : pic_data = 24'hcc3294;
          13'h0E46 : pic_data = 24'hcc328d;
          13'h0E47 : pic_data = 24'hcc327f;
          13'h0E48 : pic_data = 24'hcc3277;
          13'h0E49 : pic_data = 24'hcc3271;
          13'h0E4A : pic_data = 24'hcc3268;
          13'h0E4B : pic_data = 24'hcc3261;
          13'h0E4C : pic_data = 24'hcc3250;
          13'h0E4D : pic_data = 24'hcc3249;
          13'h0E4E : pic_data = 24'hcc3240;
          13'h0E4F : pic_data = 24'hc83536;
          13'h0E50 : pic_data = 24'hc83d36;
          13'h0E51 : pic_data = 24'hc84436;
          13'h0E52 : pic_data = 24'hc85436;
          13'h0E53 : pic_data = 24'hc85a36;
          13'h0E54 : pic_data = 24'hc86236;
          13'h0E55 : pic_data = 24'hc86936;
          13'h0E56 : pic_data = 24'hc87036;
          13'h0E57 : pic_data = 24'hc87f36;
          13'h0E58 : pic_data = 24'hc88536;
          13'h0E59 : pic_data = 24'hc88e36;
          13'h0E5A : pic_data = 24'hc89336;
          13'h0E5B : pic_data = 24'hc89b36;
          13'h0E5C : pic_data = 24'hc8ab36;
          13'h0E5D : pic_data = 24'hc8b136;
          13'h0E5E : pic_data = 24'hc8b936;
          13'h0E5F : pic_data = 24'hc8bf36;
          13'h0E60 : pic_data = 24'hcac936;
          13'h0E61 : pic_data = 24'hb9c836;
          13'h0E62 : pic_data = 24'hb3c836;
          13'h0E63 : pic_data = 24'habc836;
          13'h0E64 : pic_data = 24'h9cc836;
          13'h0E65 : pic_data = 24'h9dc836;
          13'h0E66 : pic_data = 24'h8fc836;
          13'h0E67 : pic_data = 24'h89c836;
          13'h0E68 : pic_data = 24'h80c836;
          13'h0E69 : pic_data = 24'h71c836;
          13'h0E6A : pic_data = 24'h72c836;
          13'h0E6B : pic_data = 24'h63c836;
          13'h0E6C : pic_data = 24'h5ec836;
          13'h0E6D : pic_data = 24'h53c836;
          13'h0E6E : pic_data = 24'h46c836;
          13'h0E6F : pic_data = 24'h46c836;
          13'h0E70 : pic_data = 24'h38c835;
          13'h0E71 : pic_data = 24'h35c83a;
          13'h0E72 : pic_data = 24'h36c845;
          13'h0E73 : pic_data = 24'h36c851;
          13'h0E74 : pic_data = 24'h36c858;
          13'h0E75 : pic_data = 24'h36c863;
          13'h0E76 : pic_data = 24'h36c866;
          13'h0E77 : pic_data = 24'h36c870;
          13'h0E78 : pic_data = 24'h36c87d;
          13'h0E79 : pic_data = 24'h36c883;
          13'h0E7A : pic_data = 24'h36c88e;
          13'h0E7B : pic_data = 24'h36c891;
          13'h0E7C : pic_data = 24'h36c89c;
          13'h0E7D : pic_data = 24'h36c8a7;
          13'h0E7E : pic_data = 24'h36c8af;
          13'h0E7F : pic_data = 24'h36c8ba;
          13'h0E80 : pic_data = 24'h36c8bc;
          13'h0E81 : pic_data = 24'h36caca;
          13'h0E82 : pic_data = 24'h36bdc8;
          13'h0E83 : pic_data = 24'h36b6c8;
          13'h0E84 : pic_data = 24'h36abc8;
          13'h0E85 : pic_data = 24'h369fc8;
          13'h0E86 : pic_data = 24'h369dc8;
          13'h0E87 : pic_data = 24'h3691c8;
          13'h0E88 : pic_data = 24'h368bc8;
          13'h0E89 : pic_data = 24'h3680c8;
          13'h0E8A : pic_data = 24'h3674c8;
          13'h0E8B : pic_data = 24'h3671c8;
          13'h0E8C : pic_data = 24'h3666c8;
          13'h0E8D : pic_data = 24'h3660c8;
          13'h0E8E : pic_data = 24'h3653c8;
          13'h0E8F : pic_data = 24'h3649c8;
          13'h0E90 : pic_data = 24'h3645c8;
          13'h0E91 : pic_data = 24'h363ac8;
          13'h0E92 : pic_data = 24'h3635c8;
          13'h0E93 : pic_data = 24'h4536c8;
          13'h0E94 : pic_data = 24'h4e36c8;
          13'h0E95 : pic_data = 24'h5436c8;
          13'h0E96 : pic_data = 24'h6436c8;
          13'h0E97 : pic_data = 24'h6336c8;
          13'h0E98 : pic_data = 24'h7136c8;
          13'h0E99 : pic_data = 24'h7a36c8;
          13'h0E9A : pic_data = 24'h8136c8;
          13'h0E9B : pic_data = 24'h8f36c8;
          13'h0E9C : pic_data = 24'h8d36c8;
          13'h0E9D : pic_data = 24'h9c36c8;
          13'h0E9E : pic_data = 24'ha536c8;
          13'h0E9F : pic_data = 24'hab36c8;
          13'h0EA0 : pic_data = 24'hbb36c8;
          13'h0EA1 : pic_data = 24'hb936c8;
          13'h0EA2 : pic_data = 24'hca36c9;
          13'h0EA3 : pic_data = 24'hc836bf;
          13'h0EA4 : pic_data = 24'hc836b9;
          13'h0EA5 : pic_data = 24'hc836aa;
          13'h0EA6 : pic_data = 24'hc836a3;
          13'h0EA7 : pic_data = 24'hc8369c;
          13'h0EA8 : pic_data = 24'hc83694;
          13'h0EA9 : pic_data = 24'hc8368d;
          13'h0EAA : pic_data = 24'hc8367f;
          13'h0EAB : pic_data = 24'hc83677;
          13'h0EAC : pic_data = 24'hc83671;
          13'h0EAD : pic_data = 24'hc83669;
          13'h0EAE : pic_data = 24'hc83663;
          13'h0EAF : pic_data = 24'hc83652;
          13'h0EB0 : pic_data = 24'hc8364c;
          13'h0EB1 : pic_data = 24'hc83644;
          13'h0EB2 : pic_data = 24'hc73637;
          13'h0EB3 : pic_data = 24'hc73d37;
          13'h0EB4 : pic_data = 24'hc74537;
          13'h0EB5 : pic_data = 24'hc75437;
          13'h0EB6 : pic_data = 24'hc75a37;
          13'h0EB7 : pic_data = 24'hc76337;
          13'h0EB8 : pic_data = 24'hc76a37;
          13'h0EB9 : pic_data = 24'hc77037;
          13'h0EBA : pic_data = 24'hc77f37;
          13'h0EBB : pic_data = 24'hc78537;
          13'h0EBC : pic_data = 24'hc78e37;
          13'h0EBD : pic_data = 24'hc79337;
          13'h0EBE : pic_data = 24'hc79b37;
          13'h0EBF : pic_data = 24'hc7aa37;
          13'h0EC0 : pic_data = 24'hc7b037;
          13'h0EC1 : pic_data = 24'hc7b937;
          13'h0EC2 : pic_data = 24'hc7be37;
          13'h0EC3 : pic_data = 24'hc9c937;
          13'h0EC4 : pic_data = 24'hb9c737;
          13'h0EC5 : pic_data = 24'hb3c737;
          13'h0EC6 : pic_data = 24'habc737;
          13'h0EC7 : pic_data = 24'h9cc737;
          13'h0EC8 : pic_data = 24'h9dc737;
          13'h0EC9 : pic_data = 24'h8fc737;
          13'h0ECA : pic_data = 24'h89c737;
          13'h0ECB : pic_data = 24'h80c737;
          13'h0ECC : pic_data = 24'h71c737;
          13'h0ECD : pic_data = 24'h72c737;
          13'h0ECE : pic_data = 24'h64c737;
          13'h0ECF : pic_data = 24'h5ec737;
          13'h0ED0 : pic_data = 24'h54c737;
          13'h0ED1 : pic_data = 24'h46c737;
          13'h0ED2 : pic_data = 24'h47c737;
          13'h0ED3 : pic_data = 24'h38c736;
          13'h0ED4 : pic_data = 24'h36c73b;
          13'h0ED5 : pic_data = 24'h37c745;
          13'h0ED6 : pic_data = 24'h37c751;
          13'h0ED7 : pic_data = 24'h37c758;
          13'h0ED8 : pic_data = 24'h37c763;
          13'h0ED9 : pic_data = 24'h37c766;
          13'h0EDA : pic_data = 24'h37c770;
          13'h0EDB : pic_data = 24'h37c77d;
          13'h0EDC : pic_data = 24'h37c783;
          13'h0EDD : pic_data = 24'h37c78e;
          13'h0EDE : pic_data = 24'h37c791;
          13'h0EDF : pic_data = 24'h37c79b;
          13'h0EE0 : pic_data = 24'h37c7a7;
          13'h0EE1 : pic_data = 24'h37c7ae;
          13'h0EE2 : pic_data = 24'h37c7b9;
          13'h0EE3 : pic_data = 24'h37c7bc;
          13'h0EE4 : pic_data = 24'h37c9c9;
          13'h0EE5 : pic_data = 24'h37bcc7;
          13'h0EE6 : pic_data = 24'h37b6c7;
          13'h0EE7 : pic_data = 24'h37aac7;
          13'h0EE8 : pic_data = 24'h379fc7;
          13'h0EE9 : pic_data = 24'h379cc7;
          13'h0EEA : pic_data = 24'h3791c7;
          13'h0EEB : pic_data = 24'h378bc7;
          13'h0EEC : pic_data = 24'h3780c7;
          13'h0EED : pic_data = 24'h3774c7;
          13'h0EEE : pic_data = 24'h3771c7;
          13'h0EEF : pic_data = 24'h3766c7;
          13'h0EF0 : pic_data = 24'h3760c7;
          13'h0EF1 : pic_data = 24'h3753c7;
          13'h0EF2 : pic_data = 24'h374ac7;
          13'h0EF3 : pic_data = 24'h3746c7;
          13'h0EF4 : pic_data = 24'h363bc7;
          13'h0EF5 : pic_data = 24'h3736c7;
          13'h0EF6 : pic_data = 24'h4637c7;
          13'h0EF7 : pic_data = 24'h4f37c7;
          13'h0EF8 : pic_data = 24'h5537c7;
          13'h0EF9 : pic_data = 24'h6437c7;
          13'h0EFA : pic_data = 24'h6337c7;
          13'h0EFB : pic_data = 24'h7137c7;
          13'h0EFC : pic_data = 24'h7a37c7;
          13'h0EFD : pic_data = 24'h8137c7;
          13'h0EFE : pic_data = 24'h8f37c7;
          13'h0EFF : pic_data = 24'h8d37c7;
          13'h0F00 : pic_data = 24'h9c37c7;
          13'h0F01 : pic_data = 24'ha537c7;
          13'h0F02 : pic_data = 24'hab37c7;
          13'h0F03 : pic_data = 24'hba37c7;
          13'h0F04 : pic_data = 24'hb837c7;
          13'h0F05 : pic_data = 24'hc937c9;
          13'h0F06 : pic_data = 24'hc737be;
          13'h0F07 : pic_data = 24'hc737b8;
          13'h0F08 : pic_data = 24'hc737aa;
          13'h0F09 : pic_data = 24'hc737a2;
          13'h0F0A : pic_data = 24'hc7379c;
          13'h0F0B : pic_data = 24'hc73793;
          13'h0F0C : pic_data = 24'hc7378d;
          13'h0F0D : pic_data = 24'hc7377f;
          13'h0F0E : pic_data = 24'hc73777;
          13'h0F0F : pic_data = 24'hc73771;
          13'h0F10 : pic_data = 24'hc7376a;
          13'h0F11 : pic_data = 24'hc73764;
          13'h0F12 : pic_data = 24'hc73753;
          13'h0F13 : pic_data = 24'hc7374d;
          13'h0F14 : pic_data = 24'hc73745;
          13'h0F15 : pic_data = 24'hc83536;
          13'h0F16 : pic_data = 24'hc83d36;
          13'h0F17 : pic_data = 24'hc84436;
          13'h0F18 : pic_data = 24'hc85436;
          13'h0F19 : pic_data = 24'hc85a36;
          13'h0F1A : pic_data = 24'hc86336;
          13'h0F1B : pic_data = 24'hc86936;
          13'h0F1C : pic_data = 24'hc87036;
          13'h0F1D : pic_data = 24'hc87f36;
          13'h0F1E : pic_data = 24'hc88536;
          13'h0F1F : pic_data = 24'hc88e36;
          13'h0F20 : pic_data = 24'hc89336;
          13'h0F21 : pic_data = 24'hc89b36;
          13'h0F22 : pic_data = 24'hc8ab36;
          13'h0F23 : pic_data = 24'hc8b136;
          13'h0F24 : pic_data = 24'hc8b936;
          13'h0F25 : pic_data = 24'hc8be36;
          13'h0F26 : pic_data = 24'hcac936;
          13'h0F27 : pic_data = 24'hb9c836;
          13'h0F28 : pic_data = 24'hb3c836;
          13'h0F29 : pic_data = 24'habc836;
          13'h0F2A : pic_data = 24'h9cc836;
          13'h0F2B : pic_data = 24'h9dc836;
          13'h0F2C : pic_data = 24'h8fc836;
          13'h0F2D : pic_data = 24'h89c836;
          13'h0F2E : pic_data = 24'h80c836;
          13'h0F2F : pic_data = 24'h71c836;
          13'h0F30 : pic_data = 24'h72c836;
          13'h0F31 : pic_data = 24'h64c836;
          13'h0F32 : pic_data = 24'h5ec836;
          13'h0F33 : pic_data = 24'h53c836;
          13'h0F34 : pic_data = 24'h46c836;
          13'h0F35 : pic_data = 24'h46c836;
          13'h0F36 : pic_data = 24'h38c835;
          13'h0F37 : pic_data = 24'h36c83b;
          13'h0F38 : pic_data = 24'h36c845;
          13'h0F39 : pic_data = 24'h36c851;
          13'h0F3A : pic_data = 24'h36c858;
          13'h0F3B : pic_data = 24'h36c863;
          13'h0F3C : pic_data = 24'h36c866;
          13'h0F3D : pic_data = 24'h36c870;
          13'h0F3E : pic_data = 24'h36c87d;
          13'h0F3F : pic_data = 24'h36c883;
          13'h0F40 : pic_data = 24'h36c88e;
          13'h0F41 : pic_data = 24'h36c891;
          13'h0F42 : pic_data = 24'h36c89b;
          13'h0F43 : pic_data = 24'h36c8a7;
          13'h0F44 : pic_data = 24'h36c8af;
          13'h0F45 : pic_data = 24'h36c8ba;
          13'h0F46 : pic_data = 24'h36c8bc;
          13'h0F47 : pic_data = 24'h36c9c9;
          13'h0F48 : pic_data = 24'h36bcc8;
          13'h0F49 : pic_data = 24'h36b6c8;
          13'h0F4A : pic_data = 24'h36abc8;
          13'h0F4B : pic_data = 24'h369fc8;
          13'h0F4C : pic_data = 24'h369cc8;
          13'h0F4D : pic_data = 24'h3691c8;
          13'h0F4E : pic_data = 24'h368bc8;
          13'h0F4F : pic_data = 24'h3680c8;
          13'h0F50 : pic_data = 24'h3674c8;
          13'h0F51 : pic_data = 24'h3671c8;
          13'h0F52 : pic_data = 24'h3666c8;
          13'h0F53 : pic_data = 24'h3660c8;
          13'h0F54 : pic_data = 24'h3653c8;
          13'h0F55 : pic_data = 24'h364ac8;
          13'h0F56 : pic_data = 24'h3646c8;
          13'h0F57 : pic_data = 24'h363bc8;
          13'h0F58 : pic_data = 24'h3735c8;
          13'h0F59 : pic_data = 24'h4636c8;
          13'h0F5A : pic_data = 24'h4e36c8;
          13'h0F5B : pic_data = 24'h5436c8;
          13'h0F5C : pic_data = 24'h6436c8;
          13'h0F5D : pic_data = 24'h6336c8;
          13'h0F5E : pic_data = 24'h7136c8;
          13'h0F5F : pic_data = 24'h7a36c8;
          13'h0F60 : pic_data = 24'h8136c8;
          13'h0F61 : pic_data = 24'h8f36c8;
          13'h0F62 : pic_data = 24'h8d36c8;
          13'h0F63 : pic_data = 24'h9c36c8;
          13'h0F64 : pic_data = 24'ha536c8;
          13'h0F65 : pic_data = 24'hab36c8;
          13'h0F66 : pic_data = 24'hba36c8;
          13'h0F67 : pic_data = 24'hb836c8;
          13'h0F68 : pic_data = 24'hca36c9;
          13'h0F69 : pic_data = 24'hc836bf;
          13'h0F6A : pic_data = 24'hc836b9;
          13'h0F6B : pic_data = 24'hc836aa;
          13'h0F6C : pic_data = 24'hc836a3;
          13'h0F6D : pic_data = 24'hc8369c;
          13'h0F6E : pic_data = 24'hc83693;
          13'h0F6F : pic_data = 24'hc8368d;
          13'h0F70 : pic_data = 24'hc8367f;
          13'h0F71 : pic_data = 24'hc83677;
          13'h0F72 : pic_data = 24'hc83670;
          13'h0F73 : pic_data = 24'hc83669;
          13'h0F74 : pic_data = 24'hc83663;
          13'h0F75 : pic_data = 24'hc83652;
          13'h0F76 : pic_data = 24'hc8364c;
          13'h0F77 : pic_data = 24'hc83644;
          13'h0F78 : pic_data = 24'hc43a3b;
          13'h0F79 : pic_data = 24'hc4413b;
          13'h0F7A : pic_data = 24'hc4473b;
          13'h0F7B : pic_data = 24'hc4573b;
          13'h0F7C : pic_data = 24'hc45c3b;
          13'h0F7D : pic_data = 24'hc4633b;
          13'h0F7E : pic_data = 24'hc46a3b;
          13'h0F7F : pic_data = 24'hc4713b;
          13'h0F80 : pic_data = 24'hc47f3b;
          13'h0F81 : pic_data = 24'hc4853b;
          13'h0F82 : pic_data = 24'hc48d3b;
          13'h0F83 : pic_data = 24'hc4923b;
          13'h0F84 : pic_data = 24'hc49a3b;
          13'h0F85 : pic_data = 24'hc4a83b;
          13'h0F86 : pic_data = 24'hc4ae3b;
          13'h0F87 : pic_data = 24'hc4b63b;
          13'h0F88 : pic_data = 24'hc4bc3b;
          13'h0F89 : pic_data = 24'hc6c53b;
          13'h0F8A : pic_data = 24'hb6c43b;
          13'h0F8B : pic_data = 24'hb0c43b;
          13'h0F8C : pic_data = 24'ha9c43b;
          13'h0F8D : pic_data = 24'h9bc43b;
          13'h0F8E : pic_data = 24'h9cc43b;
          13'h0F8F : pic_data = 24'h8ec43b;
          13'h0F90 : pic_data = 24'h88c43b;
          13'h0F91 : pic_data = 24'h80c43b;
          13'h0F92 : pic_data = 24'h72c43b;
          13'h0F93 : pic_data = 24'h73c43b;
          13'h0F94 : pic_data = 24'h65c43b;
          13'h0F95 : pic_data = 24'h5ec43b;
          13'h0F96 : pic_data = 24'h56c43b;
          13'h0F97 : pic_data = 24'h49c43b;
          13'h0F98 : pic_data = 24'h49c43b;
          13'h0F99 : pic_data = 24'h3cc43a;
          13'h0F9A : pic_data = 24'h3ac43e;
          13'h0F9B : pic_data = 24'h3bc448;
          13'h0F9C : pic_data = 24'h3bc453;
          13'h0F9D : pic_data = 24'h3bc45a;
          13'h0F9E : pic_data = 24'h3bc464;
          13'h0F9F : pic_data = 24'h3bc467;
          13'h0FA0 : pic_data = 24'h3bc471;
          13'h0FA1 : pic_data = 24'h3bc47d;
          13'h0FA2 : pic_data = 24'h3bc483;
          13'h0FA3 : pic_data = 24'h3bc48d;
          13'h0FA4 : pic_data = 24'h3bc490;
          13'h0FA5 : pic_data = 24'h3bc49b;
          13'h0FA6 : pic_data = 24'h3bc4a5;
          13'h0FA7 : pic_data = 24'h3bc4ac;
          13'h0FA8 : pic_data = 24'h3bc4b7;
          13'h0FA9 : pic_data = 24'h3bc4b8;
          13'h0FAA : pic_data = 24'h3bc6c6;
          13'h0FAB : pic_data = 24'h3bbac4;
          13'h0FAC : pic_data = 24'h3bb4c4;
          13'h0FAD : pic_data = 24'h3ba8c4;
          13'h0FAE : pic_data = 24'h3b9ec4;
          13'h0FAF : pic_data = 24'h3b9bc4;
          13'h0FB0 : pic_data = 24'h3b90c4;
          13'h0FB1 : pic_data = 24'h3b8ac4;
          13'h0FB2 : pic_data = 24'h3b80c4;
          13'h0FB3 : pic_data = 24'h3b75c4;
          13'h0FB4 : pic_data = 24'h3b72c4;
          13'h0FB5 : pic_data = 24'h3b67c4;
          13'h0FB6 : pic_data = 24'h3b62c4;
          13'h0FB7 : pic_data = 24'h3b56c4;
          13'h0FB8 : pic_data = 24'h3b4cc4;
          13'h0FB9 : pic_data = 24'h3b48c4;
          13'h0FBA : pic_data = 24'h3a3ec4;
          13'h0FBB : pic_data = 24'h3b3ac4;
          13'h0FBC : pic_data = 24'h483bc4;
          13'h0FBD : pic_data = 24'h513bc4;
          13'h0FBE : pic_data = 24'h573bc4;
          13'h0FBF : pic_data = 24'h643bc4;
          13'h0FC0 : pic_data = 24'h643bc4;
          13'h0FC1 : pic_data = 24'h723bc4;
          13'h0FC2 : pic_data = 24'h7b3bc4;
          13'h0FC3 : pic_data = 24'h813bc4;
          13'h0FC4 : pic_data = 24'h8e3bc4;
          13'h0FC5 : pic_data = 24'h8c3bc4;
          13'h0FC6 : pic_data = 24'h9b3bc4;
          13'h0FC7 : pic_data = 24'ha33bc4;
          13'h0FC8 : pic_data = 24'ha83bc4;
          13'h0FC9 : pic_data = 24'hb83bc4;
          13'h0FCA : pic_data = 24'hb63bc4;
          13'h0FCB : pic_data = 24'hc63bc5;
          13'h0FCC : pic_data = 24'hc43bbc;
          13'h0FCD : pic_data = 24'hc43bb6;
          13'h0FCE : pic_data = 24'hc43ba7;
          13'h0FCF : pic_data = 24'hc43ba1;
          13'h0FD0 : pic_data = 24'hc43b9b;
          13'h0FD1 : pic_data = 24'hc43b93;
          13'h0FD2 : pic_data = 24'hc43b8c;
          13'h0FD3 : pic_data = 24'hc43b7f;
          13'h0FD4 : pic_data = 24'hc43b78;
          13'h0FD5 : pic_data = 24'hc43b71;
          13'h0FD6 : pic_data = 24'hc43b6a;
          13'h0FD7 : pic_data = 24'hc43b64;
          13'h0FD8 : pic_data = 24'hc43b55;
          13'h0FD9 : pic_data = 24'hc43b4f;
          13'h0FDA : pic_data = 24'hc43b47;
          13'h0FDB : pic_data = 24'hc33b3c;
          13'h0FDC : pic_data = 24'hc3423c;
          13'h0FDD : pic_data = 24'hc3483c;
          13'h0FDE : pic_data = 24'hc3583c;
          13'h0FDF : pic_data = 24'hc35c3c;
          13'h0FE0 : pic_data = 24'hc3643c;
          13'h0FE1 : pic_data = 24'hc36b3c;
          13'h0FE2 : pic_data = 24'hc3713c;
          13'h0FE3 : pic_data = 24'hc37f3c;
          13'h0FE4 : pic_data = 24'hc3863c;
          13'h0FE5 : pic_data = 24'hc38d3c;
          13'h0FE6 : pic_data = 24'hc3923c;
          13'h0FE7 : pic_data = 24'hc39a3c;
          13'h0FE8 : pic_data = 24'hc3a73c;
          13'h0FE9 : pic_data = 24'hc3ad3c;
          13'h0FEA : pic_data = 24'hc3b63c;
          13'h0FEB : pic_data = 24'hc3bb3c;
          13'h0FEC : pic_data = 24'hc5c43c;
          13'h0FED : pic_data = 24'hb6c33c;
          13'h0FEE : pic_data = 24'hb0c33c;
          13'h0FEF : pic_data = 24'ha8c33c;
          13'h0FF0 : pic_data = 24'h9ac33c;
          13'h0FF1 : pic_data = 24'h9cc33c;
          13'h0FF2 : pic_data = 24'h8ec33c;
          13'h0FF3 : pic_data = 24'h88c33c;
          13'h0FF4 : pic_data = 24'h80c33c;
          13'h0FF5 : pic_data = 24'h72c33c;
          13'h0FF6 : pic_data = 24'h73c33c;
          13'h0FF7 : pic_data = 24'h65c33c;
          13'h0FF8 : pic_data = 24'h5fc33c;
          13'h0FF9 : pic_data = 24'h57c33c;
          13'h0FFA : pic_data = 24'h49c33c;
          13'h0FFB : pic_data = 24'h4ac33c;
          13'h0FFC : pic_data = 24'h3dc33b;
          13'h0FFD : pic_data = 24'h3bc33f;
          13'h0FFE : pic_data = 24'h3cc348;
          13'h0FFF : pic_data = 24'h3cc354;
          13'h1000 : pic_data = 24'h3cc35a;
          13'h1001 : pic_data = 24'h3cc364;
          13'h1002 : pic_data = 24'h3cc367;
          13'h1003 : pic_data = 24'h3cc371;
          13'h1004 : pic_data = 24'h3cc37d;
          13'h1005 : pic_data = 24'h3cc383;
          13'h1006 : pic_data = 24'h3cc38d;
          13'h1007 : pic_data = 24'h3cc390;
          13'h1008 : pic_data = 24'h3cc39a;
          13'h1009 : pic_data = 24'h3cc3a5;
          13'h100A : pic_data = 24'h3cc3ab;
          13'h100B : pic_data = 24'h3cc3b6;
          13'h100C : pic_data = 24'h3cc3b7;
          13'h100D : pic_data = 24'h3cc5c5;
          13'h100E : pic_data = 24'h3cb9c3;
          13'h100F : pic_data = 24'h3cb3c3;
          13'h1010 : pic_data = 24'h3ca7c3;
          13'h1011 : pic_data = 24'h3c9ec3;
          13'h1012 : pic_data = 24'h3c9bc3;
          13'h1013 : pic_data = 24'h3c90c3;
          13'h1014 : pic_data = 24'h3c8ac3;
          13'h1015 : pic_data = 24'h3c80c3;
          13'h1016 : pic_data = 24'h3c75c3;
          13'h1017 : pic_data = 24'h3c72c3;
          13'h1018 : pic_data = 24'h3c67c3;
          13'h1019 : pic_data = 24'h3c62c3;
          13'h101A : pic_data = 24'h3c56c3;
          13'h101B : pic_data = 24'h3c4dc3;
          13'h101C : pic_data = 24'h3c49c3;
          13'h101D : pic_data = 24'h3b3fc3;
          13'h101E : pic_data = 24'h3d3bc3;
          13'h101F : pic_data = 24'h493cc3;
          13'h1020 : pic_data = 24'h523cc3;
          13'h1021 : pic_data = 24'h583cc3;
          13'h1022 : pic_data = 24'h653cc3;
          13'h1023 : pic_data = 24'h643cc3;
          13'h1024 : pic_data = 24'h723cc3;
          13'h1025 : pic_data = 24'h7b3cc3;
          13'h1026 : pic_data = 24'h813cc3;
          13'h1027 : pic_data = 24'h8e3cc3;
          13'h1028 : pic_data = 24'h8c3cc3;
          13'h1029 : pic_data = 24'h9b3cc3;
          13'h102A : pic_data = 24'ha33cc3;
          13'h102B : pic_data = 24'ha83cc3;
          13'h102C : pic_data = 24'hb73cc3;
          13'h102D : pic_data = 24'hb53cc3;
          13'h102E : pic_data = 24'hc53cc4;
          13'h102F : pic_data = 24'hc33cbb;
          13'h1030 : pic_data = 24'hc33cb5;
          13'h1031 : pic_data = 24'hc33ca7;
          13'h1032 : pic_data = 24'hc33ca0;
          13'h1033 : pic_data = 24'hc33c9b;
          13'h1034 : pic_data = 24'hc33c92;
          13'h1035 : pic_data = 24'hc33c8c;
          13'h1036 : pic_data = 24'hc33c7f;
          13'h1037 : pic_data = 24'hc33c79;
          13'h1038 : pic_data = 24'hc33c72;
          13'h1039 : pic_data = 24'hc33c6b;
          13'h103A : pic_data = 24'hc33c64;
          13'h103B : pic_data = 24'hc33c56;
          13'h103C : pic_data = 24'hc33c50;
          13'h103D : pic_data = 24'hc33c48;
          13'h103E : pic_data = 24'hc43a3b;
          13'h103F : pic_data = 24'hc4413b;
          13'h1040 : pic_data = 24'hc4473b;
          13'h1041 : pic_data = 24'hc4573b;
          13'h1042 : pic_data = 24'hc45c3b;
          13'h1043 : pic_data = 24'hc4633b;
          13'h1044 : pic_data = 24'hc46a3b;
          13'h1045 : pic_data = 24'hc4713b;
          13'h1046 : pic_data = 24'hc47f3b;
          13'h1047 : pic_data = 24'hc4863b;
          13'h1048 : pic_data = 24'hc48d3b;
          13'h1049 : pic_data = 24'hc4923b;
          13'h104A : pic_data = 24'hc49a3b;
          13'h104B : pic_data = 24'hc4a73b;
          13'h104C : pic_data = 24'hc4ae3b;
          13'h104D : pic_data = 24'hc4b63b;
          13'h104E : pic_data = 24'hc4bc3b;
          13'h104F : pic_data = 24'hc6c53b;
          13'h1050 : pic_data = 24'hb6c43b;
          13'h1051 : pic_data = 24'hb0c43b;
          13'h1052 : pic_data = 24'ha8c43b;
          13'h1053 : pic_data = 24'h9ac43b;
          13'h1054 : pic_data = 24'h9cc43b;
          13'h1055 : pic_data = 24'h8ec43b;
          13'h1056 : pic_data = 24'h88c43b;
          13'h1057 : pic_data = 24'h80c43b;
          13'h1058 : pic_data = 24'h72c43b;
          13'h1059 : pic_data = 24'h73c43b;
          13'h105A : pic_data = 24'h65c43b;
          13'h105B : pic_data = 24'h5ec43b;
          13'h105C : pic_data = 24'h57c43b;
          13'h105D : pic_data = 24'h49c43b;
          13'h105E : pic_data = 24'h49c43b;
          13'h105F : pic_data = 24'h3cc43b;
          13'h1060 : pic_data = 24'h3bc43f;
          13'h1061 : pic_data = 24'h3bc448;
          13'h1062 : pic_data = 24'h3bc454;
          13'h1063 : pic_data = 24'h3bc45a;
          13'h1064 : pic_data = 24'h3bc464;
          13'h1065 : pic_data = 24'h3bc467;
          13'h1066 : pic_data = 24'h3bc471;
          13'h1067 : pic_data = 24'h3bc47d;
          13'h1068 : pic_data = 24'h3bc483;
          13'h1069 : pic_data = 24'h3bc48d;
          13'h106A : pic_data = 24'h3bc490;
          13'h106B : pic_data = 24'h3bc49b;
          13'h106C : pic_data = 24'h3bc4a5;
          13'h106D : pic_data = 24'h3bc4ab;
          13'h106E : pic_data = 24'h3bc4b7;
          13'h106F : pic_data = 24'h3bc4b8;
          13'h1070 : pic_data = 24'h3bc5c5;
          13'h1071 : pic_data = 24'h3bb9c4;
          13'h1072 : pic_data = 24'h3bb3c4;
          13'h1073 : pic_data = 24'h3ba7c4;
          13'h1074 : pic_data = 24'h3b9ec4;
          13'h1075 : pic_data = 24'h3b9bc4;
          13'h1076 : pic_data = 24'h3b90c4;
          13'h1077 : pic_data = 24'h3b8ac4;
          13'h1078 : pic_data = 24'h3b80c4;
          13'h1079 : pic_data = 24'h3b75c4;
          13'h107A : pic_data = 24'h3b72c4;
          13'h107B : pic_data = 24'h3b67c4;
          13'h107C : pic_data = 24'h3b62c4;
          13'h107D : pic_data = 24'h3b56c4;
          13'h107E : pic_data = 24'h3b4dc4;
          13'h107F : pic_data = 24'h3b49c4;
          13'h1080 : pic_data = 24'h3b3fc4;
          13'h1081 : pic_data = 24'h3c3bc4;
          13'h1082 : pic_data = 24'h483bc4;
          13'h1083 : pic_data = 24'h513bc4;
          13'h1084 : pic_data = 24'h583bc4;
          13'h1085 : pic_data = 24'h643bc4;
          13'h1086 : pic_data = 24'h643bc4;
          13'h1087 : pic_data = 24'h723bc4;
          13'h1088 : pic_data = 24'h7b3bc4;
          13'h1089 : pic_data = 24'h813bc4;
          13'h108A : pic_data = 24'h8e3bc4;
          13'h108B : pic_data = 24'h8c3bc4;
          13'h108C : pic_data = 24'h9b3bc4;
          13'h108D : pic_data = 24'ha33bc4;
          13'h108E : pic_data = 24'ha83bc4;
          13'h108F : pic_data = 24'hb73bc4;
          13'h1090 : pic_data = 24'hb53bc4;
          13'h1091 : pic_data = 24'hc63bc5;
          13'h1092 : pic_data = 24'hc43bbc;
          13'h1093 : pic_data = 24'hc43bb6;
          13'h1094 : pic_data = 24'hc43ba7;
          13'h1095 : pic_data = 24'hc43ba1;
          13'h1096 : pic_data = 24'hc43b9b;
          13'h1097 : pic_data = 24'hc43b92;
          13'h1098 : pic_data = 24'hc43b8c;
          13'h1099 : pic_data = 24'hc43b7f;
          13'h109A : pic_data = 24'hc43b79;
          13'h109B : pic_data = 24'hc43b71;
          13'h109C : pic_data = 24'hc43b6a;
          13'h109D : pic_data = 24'hc43b64;
          13'h109E : pic_data = 24'hc43b56;
          13'h109F : pic_data = 24'hc43b4f;
          13'h10A0 : pic_data = 24'hc43b47;
          13'h10A1 : pic_data = 24'hc03e3f;
          13'h10A2 : pic_data = 24'hc0453f;
          13'h10A3 : pic_data = 24'hc04b3f;
          13'h10A4 : pic_data = 24'hc0593f;
          13'h10A5 : pic_data = 24'hc05e3f;
          13'h10A6 : pic_data = 24'hc0653f;
          13'h10A7 : pic_data = 24'hc06b3f;
          13'h10A8 : pic_data = 24'hc0723f;
          13'h10A9 : pic_data = 24'hc07f3f;
          13'h10AA : pic_data = 24'hc0853f;
          13'h10AB : pic_data = 24'hc08c3f;
          13'h10AC : pic_data = 24'hc0923f;
          13'h10AD : pic_data = 24'hc0983f;
          13'h10AE : pic_data = 24'hc0a63f;
          13'h10AF : pic_data = 24'hc0ac3f;
          13'h10B0 : pic_data = 24'hc0b33f;
          13'h10B1 : pic_data = 24'hc0b83f;
          13'h10B2 : pic_data = 24'hc1c03f;
          13'h10B3 : pic_data = 24'hb3c03f;
          13'h10B4 : pic_data = 24'haec03f;
          13'h10B5 : pic_data = 24'ha6c03f;
          13'h10B6 : pic_data = 24'h99c03f;
          13'h10B7 : pic_data = 24'h9ac03f;
          13'h10B8 : pic_data = 24'h8dc03f;
          13'h10B9 : pic_data = 24'h87c03f;
          13'h10BA : pic_data = 24'h80c03f;
          13'h10BB : pic_data = 24'h73c03f;
          13'h10BC : pic_data = 24'h73c03f;
          13'h10BD : pic_data = 24'h67c03f;
          13'h10BE : pic_data = 24'h60c03f;
          13'h10BF : pic_data = 24'h58c03f;
          13'h10C0 : pic_data = 24'h4dc03f;
          13'h10C1 : pic_data = 24'h4dc03f;
          13'h10C2 : pic_data = 24'h40c03e;
          13'h10C3 : pic_data = 24'h3ec042;
          13'h10C4 : pic_data = 24'h3fc04b;
          13'h10C5 : pic_data = 24'h3fc056;
          13'h10C6 : pic_data = 24'h3fc05c;
          13'h10C7 : pic_data = 24'h3fc066;
          13'h10C8 : pic_data = 24'h3fc068;
          13'h10C9 : pic_data = 24'h3fc072;
          13'h10CA : pic_data = 24'h3fc07d;
          13'h10CB : pic_data = 24'h3fc082;
          13'h10CC : pic_data = 24'h3fc08c;
          13'h10CD : pic_data = 24'h3fc08f;
          13'h10CE : pic_data = 24'h3fc099;
          13'h10CF : pic_data = 24'h3fc0a3;
          13'h10D0 : pic_data = 24'h3fc0a9;
          13'h10D1 : pic_data = 24'h3fc0b4;
          13'h10D2 : pic_data = 24'h3fc0b5;
          13'h10D3 : pic_data = 24'h3fc1c1;
          13'h10D4 : pic_data = 24'h3fb6c0;
          13'h10D5 : pic_data = 24'h3fb1c0;
          13'h10D6 : pic_data = 24'h3fa6c0;
          13'h10D7 : pic_data = 24'h3f9cc0;
          13'h10D8 : pic_data = 24'h3f9ac0;
          13'h10D9 : pic_data = 24'h3f8fc0;
          13'h10DA : pic_data = 24'h3f8ac0;
          13'h10DB : pic_data = 24'h3f7fc0;
          13'h10DC : pic_data = 24'h3f76c0;
          13'h10DD : pic_data = 24'h3f73c0;
          13'h10DE : pic_data = 24'h3f69c0;
          13'h10DF : pic_data = 24'h3f64c0;
          13'h10E0 : pic_data = 24'h3f58c0;
          13'h10E1 : pic_data = 24'h3f4fc0;
          13'h10E2 : pic_data = 24'h3f4cc0;
          13'h10E3 : pic_data = 24'h3e42c0;
          13'h10E4 : pic_data = 24'h403ec0;
          13'h10E5 : pic_data = 24'h4c3fc0;
          13'h10E6 : pic_data = 24'h543fc0;
          13'h10E7 : pic_data = 24'h593fc0;
          13'h10E8 : pic_data = 24'h663fc0;
          13'h10E9 : pic_data = 24'h663fc0;
          13'h10EA : pic_data = 24'h733fc0;
          13'h10EB : pic_data = 24'h7b3fc0;
          13'h10EC : pic_data = 24'h803fc0;
          13'h10ED : pic_data = 24'h8d3fc0;
          13'h10EE : pic_data = 24'h8b3fc0;
          13'h10EF : pic_data = 24'h993fc0;
          13'h10F0 : pic_data = 24'ha13fc0;
          13'h10F1 : pic_data = 24'ha63fc0;
          13'h10F2 : pic_data = 24'hb53fc0;
          13'h10F3 : pic_data = 24'hb33fc0;
          13'h10F4 : pic_data = 24'hc13fc0;
          13'h10F5 : pic_data = 24'hc03fb8;
          13'h10F6 : pic_data = 24'hc03fb3;
          13'h10F7 : pic_data = 24'hc03fa5;
          13'h10F8 : pic_data = 24'hc03f9f;
          13'h10F9 : pic_data = 24'hc03f99;
          13'h10FA : pic_data = 24'hc03f92;
          13'h10FB : pic_data = 24'hc03f8c;
          13'h10FC : pic_data = 24'hc03f7f;
          13'h10FD : pic_data = 24'hc03f78;
          13'h10FE : pic_data = 24'hc03f72;
          13'h10FF : pic_data = 24'hc03f6b;
          13'h1100 : pic_data = 24'hc03f66;
          13'h1101 : pic_data = 24'hc03f57;
          13'h1102 : pic_data = 24'hc03f52;
          13'h1103 : pic_data = 24'hc03f4b;
          13'h1104 : pic_data = 24'hbe3f40;
          13'h1105 : pic_data = 24'hbe4540;
          13'h1106 : pic_data = 24'hbe4c40;
          13'h1107 : pic_data = 24'hbe5940;
          13'h1108 : pic_data = 24'hbe5e40;
          13'h1109 : pic_data = 24'hbe6640;
          13'h110A : pic_data = 24'hbe6b40;
          13'h110B : pic_data = 24'hbe7240;
          13'h110C : pic_data = 24'hbe7f40;
          13'h110D : pic_data = 24'hbe8440;
          13'h110E : pic_data = 24'hbe8c40;
          13'h110F : pic_data = 24'hbe9140;
          13'h1110 : pic_data = 24'hbe9840;
          13'h1111 : pic_data = 24'hbea540;
          13'h1112 : pic_data = 24'hbeac40;
          13'h1113 : pic_data = 24'hbeb340;
          13'h1114 : pic_data = 24'hbeb740;
          13'h1115 : pic_data = 24'hc0bf40;
          13'h1116 : pic_data = 24'hb3be40;
          13'h1117 : pic_data = 24'haebe40;
          13'h1118 : pic_data = 24'ha6be40;
          13'h1119 : pic_data = 24'h98be40;
          13'h111A : pic_data = 24'h9abe40;
          13'h111B : pic_data = 24'h8dbe40;
          13'h111C : pic_data = 24'h86be40;
          13'h111D : pic_data = 24'h80be40;
          13'h111E : pic_data = 24'h73be40;
          13'h111F : pic_data = 24'h74be40;
          13'h1120 : pic_data = 24'h67be40;
          13'h1121 : pic_data = 24'h61be40;
          13'h1122 : pic_data = 24'h59be40;
          13'h1123 : pic_data = 24'h4ebe40;
          13'h1124 : pic_data = 24'h4ebe40;
          13'h1125 : pic_data = 24'h40be3f;
          13'h1126 : pic_data = 24'h3fbe43;
          13'h1127 : pic_data = 24'h40be4c;
          13'h1128 : pic_data = 24'h40be57;
          13'h1129 : pic_data = 24'h40be5c;
          13'h112A : pic_data = 24'h40be66;
          13'h112B : pic_data = 24'h40be69;
          13'h112C : pic_data = 24'h40be72;
          13'h112D : pic_data = 24'h40be7d;
          13'h112E : pic_data = 24'h40be82;
          13'h112F : pic_data = 24'h40be8c;
          13'h1130 : pic_data = 24'h40be8f;
          13'h1131 : pic_data = 24'h40be98;
          13'h1132 : pic_data = 24'h40bea3;
          13'h1133 : pic_data = 24'h40bea8;
          13'h1134 : pic_data = 24'h40beb3;
          13'h1135 : pic_data = 24'h40beb5;
          13'h1136 : pic_data = 24'h40c0c0;
          13'h1137 : pic_data = 24'h40b5be;
          13'h1138 : pic_data = 24'h40b0be;
          13'h1139 : pic_data = 24'h40a5be;
          13'h113A : pic_data = 24'h409cbe;
          13'h113B : pic_data = 24'h4099be;
          13'h113C : pic_data = 24'h408fbe;
          13'h113D : pic_data = 24'h408abe;
          13'h113E : pic_data = 24'h407fbe;
          13'h113F : pic_data = 24'h4076be;
          13'h1140 : pic_data = 24'h4073be;
          13'h1141 : pic_data = 24'h4069be;
          13'h1142 : pic_data = 24'h4064be;
          13'h1143 : pic_data = 24'h4058be;
          13'h1144 : pic_data = 24'h4050be;
          13'h1145 : pic_data = 24'h404dbe;
          13'h1146 : pic_data = 24'h3f43be;
          13'h1147 : pic_data = 24'h403fbe;
          13'h1148 : pic_data = 24'h4d40be;
          13'h1149 : pic_data = 24'h5540be;
          13'h114A : pic_data = 24'h5a40be;
          13'h114B : pic_data = 24'h6740be;
          13'h114C : pic_data = 24'h6640be;
          13'h114D : pic_data = 24'h7340be;
          13'h114E : pic_data = 24'h7b40be;
          13'h114F : pic_data = 24'h8040be;
          13'h1150 : pic_data = 24'h8d40be;
          13'h1151 : pic_data = 24'h8b40be;
          13'h1152 : pic_data = 24'h9940be;
          13'h1153 : pic_data = 24'ha140be;
          13'h1154 : pic_data = 24'ha640be;
          13'h1155 : pic_data = 24'hb440be;
          13'h1156 : pic_data = 24'hb240be;
          13'h1157 : pic_data = 24'hc040bf;
          13'h1158 : pic_data = 24'hbe40b7;
          13'h1159 : pic_data = 24'hbe40b2;
          13'h115A : pic_data = 24'hbe40a5;
          13'h115B : pic_data = 24'hbe409e;
          13'h115C : pic_data = 24'hbe4099;
          13'h115D : pic_data = 24'hbe4091;
          13'h115E : pic_data = 24'hbe408c;
          13'h115F : pic_data = 24'hbe407f;
          13'h1160 : pic_data = 24'hbe4078;
          13'h1161 : pic_data = 24'hbe4073;
          13'h1162 : pic_data = 24'hbe406b;
          13'h1163 : pic_data = 24'hbe4066;
          13'h1164 : pic_data = 24'hbe4058;
          13'h1165 : pic_data = 24'hbe4053;
          13'h1166 : pic_data = 24'hbe404c;
          13'h1167 : pic_data = 24'hbe3f40;
          13'h1168 : pic_data = 24'hbe4640;
          13'h1169 : pic_data = 24'hbe4c40;
          13'h116A : pic_data = 24'hbe5a40;
          13'h116B : pic_data = 24'hbe5f40;
          13'h116C : pic_data = 24'hbe6640;
          13'h116D : pic_data = 24'hbe6c40;
          13'h116E : pic_data = 24'hbe7240;
          13'h116F : pic_data = 24'hbe7f40;
          13'h1170 : pic_data = 24'hbe8440;
          13'h1171 : pic_data = 24'hbe8b40;
          13'h1172 : pic_data = 24'hbe9140;
          13'h1173 : pic_data = 24'hbe9840;
          13'h1174 : pic_data = 24'hbea540;
          13'h1175 : pic_data = 24'hbeab40;
          13'h1176 : pic_data = 24'hbeb240;
          13'h1177 : pic_data = 24'hbeb740;
          13'h1178 : pic_data = 24'hbfbf40;
          13'h1179 : pic_data = 24'hb2be40;
          13'h117A : pic_data = 24'hadbe40;
          13'h117B : pic_data = 24'ha6be40;
          13'h117C : pic_data = 24'h98be40;
          13'h117D : pic_data = 24'h99be40;
          13'h117E : pic_data = 24'h8dbe40;
          13'h117F : pic_data = 24'h87be40;
          13'h1180 : pic_data = 24'h80be40;
          13'h1181 : pic_data = 24'h74be40;
          13'h1182 : pic_data = 24'h74be40;
          13'h1183 : pic_data = 24'h67be40;
          13'h1184 : pic_data = 24'h61be40;
          13'h1185 : pic_data = 24'h59be40;
          13'h1186 : pic_data = 24'h4ebe40;
          13'h1187 : pic_data = 24'h4ebe40;
          13'h1188 : pic_data = 24'h41be40;
          13'h1189 : pic_data = 24'h40be43;
          13'h118A : pic_data = 24'h40be4d;
          13'h118B : pic_data = 24'h40be57;
          13'h118C : pic_data = 24'h40be5c;
          13'h118D : pic_data = 24'h40be66;
          13'h118E : pic_data = 24'h40be69;
          13'h118F : pic_data = 24'h40be72;
          13'h1190 : pic_data = 24'h40be7d;
          13'h1191 : pic_data = 24'h40be82;
          13'h1192 : pic_data = 24'h40be8c;
          13'h1193 : pic_data = 24'h40be8f;
          13'h1194 : pic_data = 24'h40be98;
          13'h1195 : pic_data = 24'h40bea3;
          13'h1196 : pic_data = 24'h40bea8;
          13'h1197 : pic_data = 24'h40beb3;
          13'h1198 : pic_data = 24'h40beb4;
          13'h1199 : pic_data = 24'h40bfbf;
          13'h119A : pic_data = 24'h40b5be;
          13'h119B : pic_data = 24'h40afbe;
          13'h119C : pic_data = 24'h40a5be;
          13'h119D : pic_data = 24'h409cbe;
          13'h119E : pic_data = 24'h4099be;
          13'h119F : pic_data = 24'h408fbe;
          13'h11A0 : pic_data = 24'h408abe;
          13'h11A1 : pic_data = 24'h407fbe;
          13'h11A2 : pic_data = 24'h4076be;
          13'h11A3 : pic_data = 24'h4073be;
          13'h11A4 : pic_data = 24'h4069be;
          13'h11A5 : pic_data = 24'h4064be;
          13'h11A6 : pic_data = 24'h4058be;
          13'h11A7 : pic_data = 24'h4050be;
          13'h11A8 : pic_data = 24'h404ebe;
          13'h11A9 : pic_data = 24'h4043be;
          13'h11AA : pic_data = 24'h4140be;
          13'h11AB : pic_data = 24'h4d40be;
          13'h11AC : pic_data = 24'h5540be;
          13'h11AD : pic_data = 24'h5a40be;
          13'h11AE : pic_data = 24'h6740be;
          13'h11AF : pic_data = 24'h6740be;
          13'h11B0 : pic_data = 24'h7340be;
          13'h11B1 : pic_data = 24'h7b40be;
          13'h11B2 : pic_data = 24'h8040be;
          13'h11B3 : pic_data = 24'h8d40be;
          13'h11B4 : pic_data = 24'h8b40be;
          13'h11B5 : pic_data = 24'h9940be;
          13'h11B6 : pic_data = 24'ha040be;
          13'h11B7 : pic_data = 24'ha640be;
          13'h11B8 : pic_data = 24'hb340be;
          13'h11B9 : pic_data = 24'hb240be;
          13'h11BA : pic_data = 24'hbf40bf;
          13'h11BB : pic_data = 24'hbe40b7;
          13'h11BC : pic_data = 24'hbe40b2;
          13'h11BD : pic_data = 24'hbe40a5;
          13'h11BE : pic_data = 24'hbe409e;
          13'h11BF : pic_data = 24'hbe4098;
          13'h11C0 : pic_data = 24'hbe4091;
          13'h11C1 : pic_data = 24'hbe408c;
          13'h11C2 : pic_data = 24'hbe407f;
          13'h11C3 : pic_data = 24'hbe4079;
          13'h11C4 : pic_data = 24'hbe4073;
          13'h11C5 : pic_data = 24'hbe406c;
          13'h11C6 : pic_data = 24'hbe4067;
          13'h11C7 : pic_data = 24'hbe4058;
          13'h11C8 : pic_data = 24'hbe4053;
          13'h11C9 : pic_data = 24'hbe404c;
          13'h11CA : pic_data = 24'hba4344;
          13'h11CB : pic_data = 24'hba4a44;
          13'h11CC : pic_data = 24'hba4f44;
          13'h11CD : pic_data = 24'hba5b44;
          13'h11CE : pic_data = 24'hba6144;
          13'h11CF : pic_data = 24'hba6844;
          13'h11D0 : pic_data = 24'hba6e44;
          13'h11D1 : pic_data = 24'hba7344;
          13'h11D2 : pic_data = 24'hba8044;
          13'h11D3 : pic_data = 24'hba8444;
          13'h11D4 : pic_data = 24'hba8b44;
          13'h11D5 : pic_data = 24'hba8f44;
          13'h11D6 : pic_data = 24'hba9644;
          13'h11D7 : pic_data = 24'hbaa344;
          13'h11D8 : pic_data = 24'hbaa844;
          13'h11D9 : pic_data = 24'hbaae44;
          13'h11DA : pic_data = 24'hbab344;
          13'h11DB : pic_data = 24'hbbbb44;
          13'h11DC : pic_data = 24'haeba44;
          13'h11DD : pic_data = 24'haaba44;
          13'h11DE : pic_data = 24'ha4ba44;
          13'h11DF : pic_data = 24'h96ba44;
          13'h11E0 : pic_data = 24'h98ba44;
          13'h11E1 : pic_data = 24'h8bba44;
          13'h11E2 : pic_data = 24'h87ba44;
          13'h11E3 : pic_data = 24'h80ba44;
          13'h11E4 : pic_data = 24'h75ba44;
          13'h11E5 : pic_data = 24'h75ba44;
          13'h11E6 : pic_data = 24'h69ba44;
          13'h11E7 : pic_data = 24'h63ba44;
          13'h11E8 : pic_data = 24'h5bba44;
          13'h11E9 : pic_data = 24'h51ba44;
          13'h11EA : pic_data = 24'h51ba44;
          13'h11EB : pic_data = 24'h45ba43;
          13'h11EC : pic_data = 24'h44ba47;
          13'h11ED : pic_data = 24'h44ba50;
          13'h11EE : pic_data = 24'h44ba59;
          13'h11EF : pic_data = 24'h44ba5e;
          13'h11F0 : pic_data = 24'h44ba68;
          13'h11F1 : pic_data = 24'h44ba6b;
          13'h11F2 : pic_data = 24'h44ba73;
          13'h11F3 : pic_data = 24'h44ba7e;
          13'h11F4 : pic_data = 24'h44ba82;
          13'h11F5 : pic_data = 24'h44ba8b;
          13'h11F6 : pic_data = 24'h44ba8d;
          13'h11F7 : pic_data = 24'h44ba96;
          13'h11F8 : pic_data = 24'h44baa1;
          13'h11F9 : pic_data = 24'h44baa6;
          13'h11FA : pic_data = 24'h44baaf;
          13'h11FB : pic_data = 24'h44bab0;
          13'h11FC : pic_data = 24'h44bbbb;
          13'h11FD : pic_data = 24'h44b1ba;
          13'h11FE : pic_data = 24'h44abba;
          13'h11FF : pic_data = 24'h44a3ba;
          13'h1200 : pic_data = 24'h449aba;
          13'h1201 : pic_data = 24'h4497ba;
          13'h1202 : pic_data = 24'h448dba;
          13'h1203 : pic_data = 24'h4489ba;
          13'h1204 : pic_data = 24'h447fba;
          13'h1205 : pic_data = 24'h4477ba;
          13'h1206 : pic_data = 24'h4474ba;
          13'h1207 : pic_data = 24'h446bba;
          13'h1208 : pic_data = 24'h4466ba;
          13'h1209 : pic_data = 24'h445aba;
          13'h120A : pic_data = 24'h4453ba;
          13'h120B : pic_data = 24'h4450ba;
          13'h120C : pic_data = 24'h4447ba;
          13'h120D : pic_data = 24'h4543ba;
          13'h120E : pic_data = 24'h5044ba;
          13'h120F : pic_data = 24'h5744ba;
          13'h1210 : pic_data = 24'h5c44ba;
          13'h1211 : pic_data = 24'h6944ba;
          13'h1212 : pic_data = 24'h6944ba;
          13'h1213 : pic_data = 24'h7444ba;
          13'h1214 : pic_data = 24'h7b44ba;
          13'h1215 : pic_data = 24'h8044ba;
          13'h1216 : pic_data = 24'h8c44ba;
          13'h1217 : pic_data = 24'h8a44ba;
          13'h1218 : pic_data = 24'h9744ba;
          13'h1219 : pic_data = 24'h9f44ba;
          13'h121A : pic_data = 24'ha444ba;
          13'h121B : pic_data = 24'haf44ba;
          13'h121C : pic_data = 24'hae44ba;
          13'h121D : pic_data = 24'hbb44bb;
          13'h121E : pic_data = 24'hba44b3;
          13'h121F : pic_data = 24'hba44ae;
          13'h1220 : pic_data = 24'hba44a3;
          13'h1221 : pic_data = 24'hba449c;
          13'h1222 : pic_data = 24'hba4496;
          13'h1223 : pic_data = 24'hba448f;
          13'h1224 : pic_data = 24'hba448b;
          13'h1225 : pic_data = 24'hba447f;
          13'h1226 : pic_data = 24'hba447a;
          13'h1227 : pic_data = 24'hba4474;
          13'h1228 : pic_data = 24'hba446e;
          13'h1229 : pic_data = 24'hba4469;
          13'h122A : pic_data = 24'hba445a;
          13'h122B : pic_data = 24'hba4455;
          13'h122C : pic_data = 24'hba444f;
          13'h122D : pic_data = 24'hbb4343;
          13'h122E : pic_data = 24'hbb4943;
          13'h122F : pic_data = 24'hbb4f43;
          13'h1230 : pic_data = 24'hbb5b43;
          13'h1231 : pic_data = 24'hbb6043;
          13'h1232 : pic_data = 24'hbb6843;
          13'h1233 : pic_data = 24'hbb6d43;
          13'h1234 : pic_data = 24'hbb7343;
          13'h1235 : pic_data = 24'hbb8043;
          13'h1236 : pic_data = 24'hbb8443;
          13'h1237 : pic_data = 24'hbb8b43;
          13'h1238 : pic_data = 24'hbb8f43;
          13'h1239 : pic_data = 24'hbb9643;
          13'h123A : pic_data = 24'hbba343;
          13'h123B : pic_data = 24'hbba943;
          13'h123C : pic_data = 24'hbbaf43;
          13'h123D : pic_data = 24'hbbb343;
          13'h123E : pic_data = 24'hbcbb43;
          13'h123F : pic_data = 24'hafbb43;
          13'h1240 : pic_data = 24'habbb43;
          13'h1241 : pic_data = 24'ha4bb43;
          13'h1242 : pic_data = 24'h96bb43;
          13'h1243 : pic_data = 24'h98bb43;
          13'h1244 : pic_data = 24'h8bbb43;
          13'h1245 : pic_data = 24'h87bb43;
          13'h1246 : pic_data = 24'h80bb43;
          13'h1247 : pic_data = 24'h75bb43;
          13'h1248 : pic_data = 24'h74bb43;
          13'h1249 : pic_data = 24'h69bb43;
          13'h124A : pic_data = 24'h63bb43;
          13'h124B : pic_data = 24'h5bbb43;
          13'h124C : pic_data = 24'h51bb43;
          13'h124D : pic_data = 24'h50bb43;
          13'h124E : pic_data = 24'h44bb43;
          13'h124F : pic_data = 24'h43bb47;
          13'h1250 : pic_data = 24'h43bb4f;
          13'h1251 : pic_data = 24'h43bb59;
          13'h1252 : pic_data = 24'h43bb5e;
          13'h1253 : pic_data = 24'h43bb68;
          13'h1254 : pic_data = 24'h43bb6b;
          13'h1255 : pic_data = 24'h43bb73;
          13'h1256 : pic_data = 24'h43bb7e;
          13'h1257 : pic_data = 24'h43bb82;
          13'h1258 : pic_data = 24'h43bb8b;
          13'h1259 : pic_data = 24'h43bb8d;
          13'h125A : pic_data = 24'h43bb96;
          13'h125B : pic_data = 24'h43bba1;
          13'h125C : pic_data = 24'h43bba6;
          13'h125D : pic_data = 24'h43bbaf;
          13'h125E : pic_data = 24'h43bbb1;
          13'h125F : pic_data = 24'h43bcbc;
          13'h1260 : pic_data = 24'h43b1bb;
          13'h1261 : pic_data = 24'h43acbb;
          13'h1262 : pic_data = 24'h43a4bb;
          13'h1263 : pic_data = 24'h439abb;
          13'h1264 : pic_data = 24'h4397bb;
          13'h1265 : pic_data = 24'h438dbb;
          13'h1266 : pic_data = 24'h4389bb;
          13'h1267 : pic_data = 24'h437fbb;
          13'h1268 : pic_data = 24'h4377bb;
          13'h1269 : pic_data = 24'h4374bb;
          13'h126A : pic_data = 24'h436bbb;
          13'h126B : pic_data = 24'h4366bb;
          13'h126C : pic_data = 24'h435abb;
          13'h126D : pic_data = 24'h4353bb;
          13'h126E : pic_data = 24'h4350bb;
          13'h126F : pic_data = 24'h4347bb;
          13'h1270 : pic_data = 24'h4443bb;
          13'h1271 : pic_data = 24'h5043bb;
          13'h1272 : pic_data = 24'h5743bb;
          13'h1273 : pic_data = 24'h5c43bb;
          13'h1274 : pic_data = 24'h6943bb;
          13'h1275 : pic_data = 24'h6843bb;
          13'h1276 : pic_data = 24'h7443bb;
          13'h1277 : pic_data = 24'h7b43bb;
          13'h1278 : pic_data = 24'h8043bb;
          13'h1279 : pic_data = 24'h8c43bb;
          13'h127A : pic_data = 24'h8a43bb;
          13'h127B : pic_data = 24'h9743bb;
          13'h127C : pic_data = 24'h9f43bb;
          13'h127D : pic_data = 24'ha443bb;
          13'h127E : pic_data = 24'hb043bb;
          13'h127F : pic_data = 24'hae43bb;
          13'h1280 : pic_data = 24'hbc43bb;
          13'h1281 : pic_data = 24'hbb43b3;
          13'h1282 : pic_data = 24'hbb43ae;
          13'h1283 : pic_data = 24'hbb43a3;
          13'h1284 : pic_data = 24'hbb439c;
          13'h1285 : pic_data = 24'hbb4397;
          13'h1286 : pic_data = 24'hbb438f;
          13'h1287 : pic_data = 24'hbb438b;
          13'h1288 : pic_data = 24'hbb437f;
          13'h1289 : pic_data = 24'hbb437a;
          13'h128A : pic_data = 24'hbb4373;
          13'h128B : pic_data = 24'hbb436d;
          13'h128C : pic_data = 24'hbb4368;
          13'h128D : pic_data = 24'hbb435a;
          13'h128E : pic_data = 24'hbb4354;
          13'h128F : pic_data = 24'hbb434f;
          13'h1290 : pic_data = 24'hba4344;
          13'h1291 : pic_data = 24'hba4a44;
          13'h1292 : pic_data = 24'hba4f44;
          13'h1293 : pic_data = 24'hba5c44;
          13'h1294 : pic_data = 24'hba6144;
          13'h1295 : pic_data = 24'hba6844;
          13'h1296 : pic_data = 24'hba6e44;
          13'h1297 : pic_data = 24'hba7344;
          13'h1298 : pic_data = 24'hba8044;
          13'h1299 : pic_data = 24'hba8444;
          13'h129A : pic_data = 24'hba8a44;
          13'h129B : pic_data = 24'hba8f44;
          13'h129C : pic_data = 24'hba9644;
          13'h129D : pic_data = 24'hbaa344;
          13'h129E : pic_data = 24'hbaa844;
          13'h129F : pic_data = 24'hbaae44;
          13'h12A0 : pic_data = 24'hbab344;
          13'h12A1 : pic_data = 24'hbbbb44;
          13'h12A2 : pic_data = 24'haeba44;
          13'h12A3 : pic_data = 24'haaba44;
          13'h12A4 : pic_data = 24'ha4ba44;
          13'h12A5 : pic_data = 24'h96ba44;
          13'h12A6 : pic_data = 24'h98ba44;
          13'h12A7 : pic_data = 24'h8bba44;
          13'h12A8 : pic_data = 24'h87ba44;
          13'h12A9 : pic_data = 24'h80ba44;
          13'h12AA : pic_data = 24'h74ba44;
          13'h12AB : pic_data = 24'h75ba44;
          13'h12AC : pic_data = 24'h69ba44;
          13'h12AD : pic_data = 24'h63ba44;
          13'h12AE : pic_data = 24'h5bba44;
          13'h12AF : pic_data = 24'h51ba44;
          13'h12B0 : pic_data = 24'h51ba44;
          13'h12B1 : pic_data = 24'h45ba43;
          13'h12B2 : pic_data = 24'h44ba47;
          13'h12B3 : pic_data = 24'h44ba50;
          13'h12B4 : pic_data = 24'h44ba59;
          13'h12B5 : pic_data = 24'h44ba5f;
          13'h12B6 : pic_data = 24'h44ba68;
          13'h12B7 : pic_data = 24'h44ba6b;
          13'h12B8 : pic_data = 24'h44ba73;
          13'h12B9 : pic_data = 24'h44ba7e;
          13'h12BA : pic_data = 24'h44ba82;
          13'h12BB : pic_data = 24'h44ba8b;
          13'h12BC : pic_data = 24'h44ba8d;
          13'h12BD : pic_data = 24'h44ba96;
          13'h12BE : pic_data = 24'h44baa1;
          13'h12BF : pic_data = 24'h44baa6;
          13'h12C0 : pic_data = 24'h44baaf;
          13'h12C1 : pic_data = 24'h44bab0;
          13'h12C2 : pic_data = 24'h44bbbb;
          13'h12C3 : pic_data = 24'h44b1ba;
          13'h12C4 : pic_data = 24'h44abba;
          13'h12C5 : pic_data = 24'h44a3ba;
          13'h12C6 : pic_data = 24'h449aba;
          13'h12C7 : pic_data = 24'h4497ba;
          13'h12C8 : pic_data = 24'h448dba;
          13'h12C9 : pic_data = 24'h4489ba;
          13'h12CA : pic_data = 24'h447fba;
          13'h12CB : pic_data = 24'h4477ba;
          13'h12CC : pic_data = 24'h4474ba;
          13'h12CD : pic_data = 24'h446bba;
          13'h12CE : pic_data = 24'h4466ba;
          13'h12CF : pic_data = 24'h445bba;
          13'h12D0 : pic_data = 24'h4453ba;
          13'h12D1 : pic_data = 24'h4450ba;
          13'h12D2 : pic_data = 24'h4447ba;
          13'h12D3 : pic_data = 24'h4543ba;
          13'h12D4 : pic_data = 24'h5044ba;
          13'h12D5 : pic_data = 24'h5744ba;
          13'h12D6 : pic_data = 24'h5c44ba;
          13'h12D7 : pic_data = 24'h6944ba;
          13'h12D8 : pic_data = 24'h6944ba;
          13'h12D9 : pic_data = 24'h7444ba;
          13'h12DA : pic_data = 24'h7b44ba;
          13'h12DB : pic_data = 24'h8044ba;
          13'h12DC : pic_data = 24'h8b44ba;
          13'h12DD : pic_data = 24'h8a44ba;
          13'h12DE : pic_data = 24'h9744ba;
          13'h12DF : pic_data = 24'h9e44ba;
          13'h12E0 : pic_data = 24'ha344ba;
          13'h12E1 : pic_data = 24'haf44ba;
          13'h12E2 : pic_data = 24'hae44ba;
          13'h12E3 : pic_data = 24'hbb44bb;
          13'h12E4 : pic_data = 24'hba44b3;
          13'h12E5 : pic_data = 24'hba44ae;
          13'h12E6 : pic_data = 24'hba44a3;
          13'h12E7 : pic_data = 24'hba449c;
          13'h12E8 : pic_data = 24'hba4497;
          13'h12E9 : pic_data = 24'hba448f;
          13'h12EA : pic_data = 24'hba448b;
          13'h12EB : pic_data = 24'hba447f;
          13'h12EC : pic_data = 24'hba4479;
          13'h12ED : pic_data = 24'hba4474;
          13'h12EE : pic_data = 24'hba446e;
          13'h12EF : pic_data = 24'hba4468;
          13'h12F0 : pic_data = 24'hba445a;
          13'h12F1 : pic_data = 24'hba4455;
          13'h12F2 : pic_data = 24'hba444f;
          13'h12F3 : pic_data = 24'hb64748;
          13'h12F4 : pic_data = 24'hb64d48;
          13'h12F5 : pic_data = 24'hb65248;
          13'h12F6 : pic_data = 24'hb66048;
          13'h12F7 : pic_data = 24'hb66448;
          13'h12F8 : pic_data = 24'hb66848;
          13'h12F9 : pic_data = 24'hb66f48;
          13'h12FA : pic_data = 24'hb67448;
          13'h12FB : pic_data = 24'hb68048;
          13'h12FC : pic_data = 24'hb68548;
          13'h12FD : pic_data = 24'hb68948;
          13'h12FE : pic_data = 24'hb68e48;
          13'h12FF : pic_data = 24'hb69548;
          13'h1300 : pic_data = 24'hb69e48;
          13'h1301 : pic_data = 24'hb6a448;
          13'h1302 : pic_data = 24'hb6ab48;
          13'h1303 : pic_data = 24'hb6b048;
          13'h1304 : pic_data = 24'hb7b748;
          13'h1305 : pic_data = 24'hacb648;
          13'h1306 : pic_data = 24'ha6b648;
          13'h1307 : pic_data = 24'h9fb648;
          13'h1308 : pic_data = 24'h95b648;
          13'h1309 : pic_data = 24'h97b648;
          13'h130A : pic_data = 24'h8ab648;
          13'h130B : pic_data = 24'h86b648;
          13'h130C : pic_data = 24'h80b648;
          13'h130D : pic_data = 24'h74b648;
          13'h130E : pic_data = 24'h76b648;
          13'h130F : pic_data = 24'h6ab648;
          13'h1310 : pic_data = 24'h65b648;
          13'h1311 : pic_data = 24'h5fb648;
          13'h1312 : pic_data = 24'h54b648;
          13'h1313 : pic_data = 24'h54b648;
          13'h1314 : pic_data = 24'h49b647;
          13'h1315 : pic_data = 24'h48b64c;
          13'h1316 : pic_data = 24'h48b652;
          13'h1317 : pic_data = 24'h48b65e;
          13'h1318 : pic_data = 24'h48b662;
          13'h1319 : pic_data = 24'h48b669;
          13'h131A : pic_data = 24'h48b66c;
          13'h131B : pic_data = 24'h48b674;
          13'h131C : pic_data = 24'h48b67e;
          13'h131D : pic_data = 24'h48b682;
          13'h131E : pic_data = 24'h48b68a;
          13'h131F : pic_data = 24'h48b68c;
          13'h1320 : pic_data = 24'h48b696;
          13'h1321 : pic_data = 24'h48b69e;
          13'h1322 : pic_data = 24'h48b6a2;
          13'h1323 : pic_data = 24'h48b6ac;
          13'h1324 : pic_data = 24'h48b6ae;
          13'h1325 : pic_data = 24'h48b7b7;
          13'h1326 : pic_data = 24'h48aeb6;
          13'h1327 : pic_data = 24'h48a9b6;
          13'h1328 : pic_data = 24'h489fb6;
          13'h1329 : pic_data = 24'h4898b6;
          13'h132A : pic_data = 24'h4896b6;
          13'h132B : pic_data = 24'h488cb6;
          13'h132C : pic_data = 24'h4888b6;
          13'h132D : pic_data = 24'h4880b6;
          13'h132E : pic_data = 24'h4877b6;
          13'h132F : pic_data = 24'h4875b6;
          13'h1330 : pic_data = 24'h486cb6;
          13'h1331 : pic_data = 24'h4867b6;
          13'h1332 : pic_data = 24'h485fb6;
          13'h1333 : pic_data = 24'h4856b6;
          13'h1334 : pic_data = 24'h4853b6;
          13'h1335 : pic_data = 24'h484cb6;
          13'h1336 : pic_data = 24'h4947b6;
          13'h1337 : pic_data = 24'h5348b6;
          13'h1338 : pic_data = 24'h5b48b6;
          13'h1339 : pic_data = 24'h5f48b6;
          13'h133A : pic_data = 24'h6948b6;
          13'h133B : pic_data = 24'h6a48b6;
          13'h133C : pic_data = 24'h7548b6;
          13'h133D : pic_data = 24'h7c48b6;
          13'h133E : pic_data = 24'h8048b6;
          13'h133F : pic_data = 24'h8a48b6;
          13'h1340 : pic_data = 24'h8948b6;
          13'h1341 : pic_data = 24'h9648b6;
          13'h1342 : pic_data = 24'h9b48b6;
          13'h1343 : pic_data = 24'h9f48b6;
          13'h1344 : pic_data = 24'hac48b6;
          13'h1345 : pic_data = 24'hab48b6;
          13'h1346 : pic_data = 24'hb748b7;
          13'h1347 : pic_data = 24'hb648b0;
          13'h1348 : pic_data = 24'hb648ab;
          13'h1349 : pic_data = 24'hb6489e;
          13'h134A : pic_data = 24'hb64899;
          13'h134B : pic_data = 24'hb64896;
          13'h134C : pic_data = 24'hb6488e;
          13'h134D : pic_data = 24'hb6488a;
          13'h134E : pic_data = 24'hb6487f;
          13'h134F : pic_data = 24'hb64879;
          13'h1350 : pic_data = 24'hb64875;
          13'h1351 : pic_data = 24'hb6486f;
          13'h1352 : pic_data = 24'hb64869;
          13'h1353 : pic_data = 24'hb6485e;
          13'h1354 : pic_data = 24'hb64859;
          13'h1355 : pic_data = 24'hb64852;
          13'h1356 : pic_data = 24'hb74747;
          13'h1357 : pic_data = 24'hb74c47;
          13'h1358 : pic_data = 24'hb75247;
          13'h1359 : pic_data = 24'hb75f47;
          13'h135A : pic_data = 24'hb76347;
          13'h135B : pic_data = 24'hb76847;
          13'h135C : pic_data = 24'hb76e47;
          13'h135D : pic_data = 24'hb77447;
          13'h135E : pic_data = 24'hb78047;
          13'h135F : pic_data = 24'hb78547;
          13'h1360 : pic_data = 24'hb78a47;
          13'h1361 : pic_data = 24'hb78e47;
          13'h1362 : pic_data = 24'hb79547;
          13'h1363 : pic_data = 24'hb79f47;
          13'h1364 : pic_data = 24'hb7a447;
          13'h1365 : pic_data = 24'hb7ac47;
          13'h1366 : pic_data = 24'hb7b047;
          13'h1367 : pic_data = 24'hb8b747;
          13'h1368 : pic_data = 24'hacb747;
          13'h1369 : pic_data = 24'ha7b747;
          13'h136A : pic_data = 24'ha0b747;
          13'h136B : pic_data = 24'h96b747;
          13'h136C : pic_data = 24'h97b747;
          13'h136D : pic_data = 24'h8ab747;
          13'h136E : pic_data = 24'h86b747;
          13'h136F : pic_data = 24'h80b747;
          13'h1370 : pic_data = 24'h74b747;
          13'h1371 : pic_data = 24'h76b747;
          13'h1372 : pic_data = 24'h6ab747;
          13'h1373 : pic_data = 24'h64b747;
          13'h1374 : pic_data = 24'h5fb747;
          13'h1375 : pic_data = 24'h53b747;
          13'h1376 : pic_data = 24'h53b747;
          13'h1377 : pic_data = 24'h49b747;
          13'h1378 : pic_data = 24'h47b74b;
          13'h1379 : pic_data = 24'h47b752;
          13'h137A : pic_data = 24'h47b75d;
          13'h137B : pic_data = 24'h47b761;
          13'h137C : pic_data = 24'h47b769;
          13'h137D : pic_data = 24'h47b76c;
          13'h137E : pic_data = 24'h47b774;
          13'h137F : pic_data = 24'h47b77e;
          13'h1380 : pic_data = 24'h47b782;
          13'h1381 : pic_data = 24'h47b78a;
          13'h1382 : pic_data = 24'h47b78c;
          13'h1383 : pic_data = 24'h47b796;
          13'h1384 : pic_data = 24'h47b79e;
          13'h1385 : pic_data = 24'h47b7a2;
          13'h1386 : pic_data = 24'h47b7ac;
          13'h1387 : pic_data = 24'h47b7ae;
          13'h1388 : pic_data = 24'h47b8b8;
          13'h1389 : pic_data = 24'h47aeb7;
          13'h138A : pic_data = 24'h47a9b7;
          13'h138B : pic_data = 24'h479fb7;
          13'h138C : pic_data = 24'h4798b7;
          13'h138D : pic_data = 24'h4796b7;
          13'h138E : pic_data = 24'h478cb7;
          13'h138F : pic_data = 24'h4788b7;
          13'h1390 : pic_data = 24'h4780b7;
          13'h1391 : pic_data = 24'h4777b7;
          13'h1392 : pic_data = 24'h4775b7;
          13'h1393 : pic_data = 24'h476cb7;
          13'h1394 : pic_data = 24'h4767b7;
          13'h1395 : pic_data = 24'h475eb7;
          13'h1396 : pic_data = 24'h4756b7;
          13'h1397 : pic_data = 24'h4753b7;
          13'h1398 : pic_data = 24'h474bb7;
          13'h1399 : pic_data = 24'h4947b7;
          13'h139A : pic_data = 24'h5347b7;
          13'h139B : pic_data = 24'h5b47b7;
          13'h139C : pic_data = 24'h5f47b7;
          13'h139D : pic_data = 24'h6947b7;
          13'h139E : pic_data = 24'h6947b7;
          13'h139F : pic_data = 24'h7547b7;
          13'h13A0 : pic_data = 24'h7c47b7;
          13'h13A1 : pic_data = 24'h8047b7;
          13'h13A2 : pic_data = 24'h8b47b7;
          13'h13A3 : pic_data = 24'h8947b7;
          13'h13A4 : pic_data = 24'h9647b7;
          13'h13A5 : pic_data = 24'h9c47b7;
          13'h13A6 : pic_data = 24'ha047b7;
          13'h13A7 : pic_data = 24'had47b7;
          13'h13A8 : pic_data = 24'hab47b7;
          13'h13A9 : pic_data = 24'hb847b7;
          13'h13AA : pic_data = 24'hb747b1;
          13'h13AB : pic_data = 24'hb747ab;
          13'h13AC : pic_data = 24'hb7479f;
          13'h13AD : pic_data = 24'hb74799;
          13'h13AE : pic_data = 24'hb74796;
          13'h13AF : pic_data = 24'hb7478e;
          13'h13B0 : pic_data = 24'hb7478a;
          13'h13B1 : pic_data = 24'hb7477f;
          13'h13B2 : pic_data = 24'hb74779;
          13'h13B3 : pic_data = 24'hb74775;
          13'h13B4 : pic_data = 24'hb7476e;
          13'h13B5 : pic_data = 24'hb74769;
          13'h13B6 : pic_data = 24'hb7475e;
          13'h13B7 : pic_data = 24'hb74758;
          13'h13B8 : pic_data = 24'hb74752;
          13'h13B9 : pic_data = 24'hb64748;
          13'h13BA : pic_data = 24'hb64d48;
          13'h13BB : pic_data = 24'hb65248;
          13'h13BC : pic_data = 24'hb66048;
          13'h13BD : pic_data = 24'hb66448;
          13'h13BE : pic_data = 24'hb66948;
          13'h13BF : pic_data = 24'hb66f48;
          13'h13C0 : pic_data = 24'hb67448;
          13'h13C1 : pic_data = 24'hb68048;
          13'h13C2 : pic_data = 24'hb68548;
          13'h13C3 : pic_data = 24'hb68a48;
          13'h13C4 : pic_data = 24'hb68e48;
          13'h13C5 : pic_data = 24'hb69548;
          13'h13C6 : pic_data = 24'hb69f48;
          13'h13C7 : pic_data = 24'hb6a448;
          13'h13C8 : pic_data = 24'hb6ab48;
          13'h13C9 : pic_data = 24'hb6b048;
          13'h13CA : pic_data = 24'hb7b748;
          13'h13CB : pic_data = 24'hacb648;
          13'h13CC : pic_data = 24'ha6b648;
          13'h13CD : pic_data = 24'ha0b648;
          13'h13CE : pic_data = 24'h95b648;
          13'h13CF : pic_data = 24'h97b648;
          13'h13D0 : pic_data = 24'h8ab648;
          13'h13D1 : pic_data = 24'h86b648;
          13'h13D2 : pic_data = 24'h80b648;
          13'h13D3 : pic_data = 24'h74b648;
          13'h13D4 : pic_data = 24'h76b648;
          13'h13D5 : pic_data = 24'h6ab648;
          13'h13D6 : pic_data = 24'h65b648;
          13'h13D7 : pic_data = 24'h5fb648;
          13'h13D8 : pic_data = 24'h54b648;
          13'h13D9 : pic_data = 24'h54b648;
          13'h13DA : pic_data = 24'h49b647;
          13'h13DB : pic_data = 24'h48b64b;
          13'h13DC : pic_data = 24'h48b653;
          13'h13DD : pic_data = 24'h48b65d;
          13'h13DE : pic_data = 24'h48b661;
          13'h13DF : pic_data = 24'h48b669;
          13'h13E0 : pic_data = 24'h48b66c;
          13'h13E1 : pic_data = 24'h48b674;
          13'h13E2 : pic_data = 24'h48b67e;
          13'h13E3 : pic_data = 24'h48b682;
          13'h13E4 : pic_data = 24'h48b68a;
          13'h13E5 : pic_data = 24'h48b68c;
          13'h13E6 : pic_data = 24'h48b695;
          13'h13E7 : pic_data = 24'h48b69e;
          13'h13E8 : pic_data = 24'h48b6a2;
          13'h13E9 : pic_data = 24'h48b6ac;
          13'h13EA : pic_data = 24'h48b6ad;
          13'h13EB : pic_data = 24'h48b7b7;
          13'h13EC : pic_data = 24'h48aeb6;
          13'h13ED : pic_data = 24'h48a9b6;
          13'h13EE : pic_data = 24'h489fb6;
          13'h13EF : pic_data = 24'h4898b6;
          13'h13F0 : pic_data = 24'h4896b6;
          13'h13F1 : pic_data = 24'h488cb6;
          13'h13F2 : pic_data = 24'h4888b6;
          13'h13F3 : pic_data = 24'h4880b6;
          13'h13F4 : pic_data = 24'h4877b6;
          13'h13F5 : pic_data = 24'h4875b6;
          13'h13F6 : pic_data = 24'h486cb6;
          13'h13F7 : pic_data = 24'h4867b6;
          13'h13F8 : pic_data = 24'h485fb6;
          13'h13F9 : pic_data = 24'h4856b6;
          13'h13FA : pic_data = 24'h4853b6;
          13'h13FB : pic_data = 24'h484bb6;
          13'h13FC : pic_data = 24'h4947b6;
          13'h13FD : pic_data = 24'h5348b6;
          13'h13FE : pic_data = 24'h5b48b6;
          13'h13FF : pic_data = 24'h5f48b6;
          13'h1400 : pic_data = 24'h6a48b6;
          13'h1401 : pic_data = 24'h6a48b6;
          13'h1402 : pic_data = 24'h7548b6;
          13'h1403 : pic_data = 24'h7c48b6;
          13'h1404 : pic_data = 24'h8048b6;
          13'h1405 : pic_data = 24'h8b48b6;
          13'h1406 : pic_data = 24'h8948b6;
          13'h1407 : pic_data = 24'h9648b6;
          13'h1408 : pic_data = 24'h9b48b6;
          13'h1409 : pic_data = 24'ha048b6;
          13'h140A : pic_data = 24'hac48b6;
          13'h140B : pic_data = 24'hab48b6;
          13'h140C : pic_data = 24'hb748b7;
          13'h140D : pic_data = 24'hb648b0;
          13'h140E : pic_data = 24'hb648ab;
          13'h140F : pic_data = 24'hb6489f;
          13'h1410 : pic_data = 24'hb64899;
          13'h1411 : pic_data = 24'hb64896;
          13'h1412 : pic_data = 24'hb6488e;
          13'h1413 : pic_data = 24'hb6488a;
          13'h1414 : pic_data = 24'hb6487f;
          13'h1415 : pic_data = 24'hb64879;
          13'h1416 : pic_data = 24'hb64875;
          13'h1417 : pic_data = 24'hb6486f;
          13'h1418 : pic_data = 24'hb64869;
          13'h1419 : pic_data = 24'hb6485e;
          13'h141A : pic_data = 24'hb64859;
          13'h141B : pic_data = 24'hb64852;
          13'h141C : pic_data = 24'hb24c4d;
          13'h141D : pic_data = 24'hb2524d;
          13'h141E : pic_data = 24'hb2564d;
          13'h141F : pic_data = 24'hb2614d;
          13'h1420 : pic_data = 24'hb2664d;
          13'h1421 : pic_data = 24'hb26b4d;
          13'h1422 : pic_data = 24'hb2704d;
          13'h1423 : pic_data = 24'hb2744d;
          13'h1424 : pic_data = 24'hb2804d;
          13'h1425 : pic_data = 24'hb2854d;
          13'h1426 : pic_data = 24'hb28a4d;
          13'h1427 : pic_data = 24'hb28d4d;
          13'h1428 : pic_data = 24'hb2934d;
          13'h1429 : pic_data = 24'hb29d4d;
          13'h142A : pic_data = 24'hb2a14d;
          13'h142B : pic_data = 24'hb2a74d;
          13'h142C : pic_data = 24'hb2ac4d;
          13'h142D : pic_data = 24'hb3b34d;
          13'h142E : pic_data = 24'ha7b24d;
          13'h142F : pic_data = 24'ha3b24d;
          13'h1430 : pic_data = 24'h9eb24d;
          13'h1431 : pic_data = 24'h93b24d;
          13'h1432 : pic_data = 24'h94b24d;
          13'h1433 : pic_data = 24'h8ab24d;
          13'h1434 : pic_data = 24'h86b24d;
          13'h1435 : pic_data = 24'h80b24d;
          13'h1436 : pic_data = 24'h74b24d;
          13'h1437 : pic_data = 24'h76b24d;
          13'h1438 : pic_data = 24'h6bb24d;
          13'h1439 : pic_data = 24'h67b24d;
          13'h143A : pic_data = 24'h61b24d;
          13'h143B : pic_data = 24'h58b24d;
          13'h143C : pic_data = 24'h58b24d;
          13'h143D : pic_data = 24'h4eb24d;
          13'h143E : pic_data = 24'h4db24f;
          13'h143F : pic_data = 24'h4db257;
          13'h1440 : pic_data = 24'h4db25f;
          13'h1441 : pic_data = 24'h4db263;
          13'h1442 : pic_data = 24'h4db26b;
          13'h1443 : pic_data = 24'h4db26d;
          13'h1444 : pic_data = 24'h4db274;
          13'h1445 : pic_data = 24'h4db27e;
          13'h1446 : pic_data = 24'h4db282;
          13'h1447 : pic_data = 24'h4db28a;
          13'h1448 : pic_data = 24'h4db28c;
          13'h1449 : pic_data = 24'h4db293;
          13'h144A : pic_data = 24'h4db29c;
          13'h144B : pic_data = 24'h4db2a0;
          13'h144C : pic_data = 24'h4db2a8;
          13'h144D : pic_data = 24'h4db2a9;
          13'h144E : pic_data = 24'h4db3b3;
          13'h144F : pic_data = 24'h4daab2;
          13'h1450 : pic_data = 24'h4da6b2;
          13'h1451 : pic_data = 24'h4d9db2;
          13'h1452 : pic_data = 24'h4d96b2;
          13'h1453 : pic_data = 24'h4d94b2;
          13'h1454 : pic_data = 24'h4d8cb2;
          13'h1455 : pic_data = 24'h4d88b2;
          13'h1456 : pic_data = 24'h4d80b2;
          13'h1457 : pic_data = 24'h4d77b2;
          13'h1458 : pic_data = 24'h4d75b2;
          13'h1459 : pic_data = 24'h4d6db2;
          13'h145A : pic_data = 24'h4d69b2;
          13'h145B : pic_data = 24'h4d61b2;
          13'h145C : pic_data = 24'h4d59b2;
          13'h145D : pic_data = 24'h4d57b2;
          13'h145E : pic_data = 24'h4d4fb2;
          13'h145F : pic_data = 24'h4e4db2;
          13'h1460 : pic_data = 24'h574db2;
          13'h1461 : pic_data = 24'h5d4db2;
          13'h1462 : pic_data = 24'h614db2;
          13'h1463 : pic_data = 24'h6c4db2;
          13'h1464 : pic_data = 24'h6b4db2;
          13'h1465 : pic_data = 24'h754db2;
          13'h1466 : pic_data = 24'h7c4db2;
          13'h1467 : pic_data = 24'h804db2;
          13'h1468 : pic_data = 24'h8b4db2;
          13'h1469 : pic_data = 24'h8a4db2;
          13'h146A : pic_data = 24'h944db2;
          13'h146B : pic_data = 24'h994db2;
          13'h146C : pic_data = 24'h9e4db2;
          13'h146D : pic_data = 24'ha84db2;
          13'h146E : pic_data = 24'ha74db2;
          13'h146F : pic_data = 24'hb34db3;
          13'h1470 : pic_data = 24'hb24dac;
          13'h1471 : pic_data = 24'hb24da6;
          13'h1472 : pic_data = 24'hb24d9d;
          13'h1473 : pic_data = 24'hb24d97;
          13'h1474 : pic_data = 24'hb24d93;
          13'h1475 : pic_data = 24'hb24d8f;
          13'h1476 : pic_data = 24'hb24d8a;
          13'h1477 : pic_data = 24'hb24d7f;
          13'h1478 : pic_data = 24'hb24d79;
          13'h1479 : pic_data = 24'hb24d75;
          13'h147A : pic_data = 24'hb24d70;
          13'h147B : pic_data = 24'hb24d6b;
          13'h147C : pic_data = 24'hb24d60;
          13'h147D : pic_data = 24'hb24d5c;
          13'h147E : pic_data = 24'hb24d56;
          13'h147F : pic_data = 24'hb34c4c;
          13'h1480 : pic_data = 24'hb3514c;
          13'h1481 : pic_data = 24'hb3564c;
          13'h1482 : pic_data = 24'hb3614c;
          13'h1483 : pic_data = 24'hb3654c;
          13'h1484 : pic_data = 24'hb36a4c;
          13'h1485 : pic_data = 24'hb36f4c;
          13'h1486 : pic_data = 24'hb3744c;
          13'h1487 : pic_data = 24'hb3804c;
          13'h1488 : pic_data = 24'hb3854c;
          13'h1489 : pic_data = 24'hb38a4c;
          13'h148A : pic_data = 24'hb38d4c;
          13'h148B : pic_data = 24'hb3934c;
          13'h148C : pic_data = 24'hb39d4c;
          13'h148D : pic_data = 24'hb3a24c;
          13'h148E : pic_data = 24'hb3a84c;
          13'h148F : pic_data = 24'hb3ad4c;
          13'h1490 : pic_data = 24'hb4b44c;
          13'h1491 : pic_data = 24'ha8b34c;
          13'h1492 : pic_data = 24'ha4b34c;
          13'h1493 : pic_data = 24'h9eb34c;
          13'h1494 : pic_data = 24'h94b34c;
          13'h1495 : pic_data = 24'h95b34c;
          13'h1496 : pic_data = 24'h8ab34c;
          13'h1497 : pic_data = 24'h86b34c;
          13'h1498 : pic_data = 24'h80b34c;
          13'h1499 : pic_data = 24'h74b34c;
          13'h149A : pic_data = 24'h75b34c;
          13'h149B : pic_data = 24'h6bb34c;
          13'h149C : pic_data = 24'h66b34c;
          13'h149D : pic_data = 24'h61b34c;
          13'h149E : pic_data = 24'h58b34c;
          13'h149F : pic_data = 24'h57b34c;
          13'h14A0 : pic_data = 24'h4db34c;
          13'h14A1 : pic_data = 24'h4cb34f;
          13'h14A2 : pic_data = 24'h4cb356;
          13'h14A3 : pic_data = 24'h4cb35f;
          13'h14A4 : pic_data = 24'h4cb363;
          13'h14A5 : pic_data = 24'h4cb36b;
          13'h14A6 : pic_data = 24'h4cb36d;
          13'h14A7 : pic_data = 24'h4cb374;
          13'h14A8 : pic_data = 24'h4cb37e;
          13'h14A9 : pic_data = 24'h4cb382;
          13'h14AA : pic_data = 24'h4cb38a;
          13'h14AB : pic_data = 24'h4cb38c;
          13'h14AC : pic_data = 24'h4cb393;
          13'h14AD : pic_data = 24'h4cb39c;
          13'h14AE : pic_data = 24'h4cb3a0;
          13'h14AF : pic_data = 24'h4cb3a8;
          13'h14B0 : pic_data = 24'h4cb3aa;
          13'h14B1 : pic_data = 24'h4cb4b4;
          13'h14B2 : pic_data = 24'h4caab3;
          13'h14B3 : pic_data = 24'h4ca6b3;
          13'h14B4 : pic_data = 24'h4c9eb3;
          13'h14B5 : pic_data = 24'h4c96b3;
          13'h14B6 : pic_data = 24'h4c94b3;
          13'h14B7 : pic_data = 24'h4c8cb3;
          13'h14B8 : pic_data = 24'h4c88b3;
          13'h14B9 : pic_data = 24'h4c80b3;
          13'h14BA : pic_data = 24'h4c77b3;
          13'h14BB : pic_data = 24'h4c75b3;
          13'h14BC : pic_data = 24'h4c6db3;
          13'h14BD : pic_data = 24'h4c69b3;
          13'h14BE : pic_data = 24'h4c60b3;
          13'h14BF : pic_data = 24'h4c59b3;
          13'h14C0 : pic_data = 24'h4c57b3;
          13'h14C1 : pic_data = 24'h4c4fb3;
          13'h14C2 : pic_data = 24'h4e4cb3;
          13'h14C3 : pic_data = 24'h574cb3;
          13'h14C4 : pic_data = 24'h5c4cb3;
          13'h14C5 : pic_data = 24'h614cb3;
          13'h14C6 : pic_data = 24'h6b4cb3;
          13'h14C7 : pic_data = 24'h6a4cb3;
          13'h14C8 : pic_data = 24'h754cb3;
          13'h14C9 : pic_data = 24'h7c4cb3;
          13'h14CA : pic_data = 24'h804cb3;
          13'h14CB : pic_data = 24'h8b4cb3;
          13'h14CC : pic_data = 24'h8a4cb3;
          13'h14CD : pic_data = 24'h944cb3;
          13'h14CE : pic_data = 24'h9a4cb3;
          13'h14CF : pic_data = 24'h9e4cb3;
          13'h14D0 : pic_data = 24'ha94cb3;
          13'h14D1 : pic_data = 24'ha84cb3;
          13'h14D2 : pic_data = 24'hb44cb4;
          13'h14D3 : pic_data = 24'hb34cad;
          13'h14D4 : pic_data = 24'hb34ca7;
          13'h14D5 : pic_data = 24'hb34c9d;
          13'h14D6 : pic_data = 24'hb34c97;
          13'h14D7 : pic_data = 24'hb34c94;
          13'h14D8 : pic_data = 24'hb34c8f;
          13'h14D9 : pic_data = 24'hb34c8a;
          13'h14DA : pic_data = 24'hb34c7f;
          13'h14DB : pic_data = 24'hb34c79;
          13'h14DC : pic_data = 24'hb34c74;
          13'h14DD : pic_data = 24'hb34c6f;
          13'h14DE : pic_data = 24'hb34c6b;
          13'h14DF : pic_data = 24'hb34c60;
          13'h14E0 : pic_data = 24'hb34c5b;
          13'h14E1 : pic_data = 24'hb34c56;
          13'h14E2 : pic_data = 24'haf4f4f;
          13'h14E3 : pic_data = 24'haf544f;
          13'h14E4 : pic_data = 24'haf584f;
          13'h14E5 : pic_data = 24'haf634f;
          13'h14E6 : pic_data = 24'haf674f;
          13'h14E7 : pic_data = 24'haf6b4f;
          13'h14E8 : pic_data = 24'haf704f;
          13'h14E9 : pic_data = 24'haf754f;
          13'h14EA : pic_data = 24'haf804f;
          13'h14EB : pic_data = 24'haf844f;
          13'h14EC : pic_data = 24'haf894f;
          13'h14ED : pic_data = 24'haf8d4f;
          13'h14EE : pic_data = 24'haf934f;
          13'h14EF : pic_data = 24'haf9b4f;
          13'h14F0 : pic_data = 24'haf9f4f;
          13'h14F1 : pic_data = 24'hafa64f;
          13'h14F2 : pic_data = 24'hafaa4f;
          13'h14F3 : pic_data = 24'hb0b04f;
          13'h14F4 : pic_data = 24'ha6af4f;
          13'h14F5 : pic_data = 24'ha2af4f;
          13'h14F6 : pic_data = 24'h9caf4f;
          13'h14F7 : pic_data = 24'h93af4f;
          13'h14F8 : pic_data = 24'h94af4f;
          13'h14F9 : pic_data = 24'h89af4f;
          13'h14FA : pic_data = 24'h86af4f;
          13'h14FB : pic_data = 24'h80af4f;
          13'h14FC : pic_data = 24'h75af4f;
          13'h14FD : pic_data = 24'h76af4f;
          13'h14FE : pic_data = 24'h6caf4f;
          13'h14FF : pic_data = 24'h68af4f;
          13'h1500 : pic_data = 24'h63af4f;
          13'h1501 : pic_data = 24'h5aaf4f;
          13'h1502 : pic_data = 24'h59af4f;
          13'h1503 : pic_data = 24'h51af4f;
          13'h1504 : pic_data = 24'h4faf52;
          13'h1505 : pic_data = 24'h4faf58;
          13'h1506 : pic_data = 24'h4faf61;
          13'h1507 : pic_data = 24'h4faf65;
          13'h1508 : pic_data = 24'h4faf6c;
          13'h1509 : pic_data = 24'h4faf6e;
          13'h150A : pic_data = 24'h4faf75;
          13'h150B : pic_data = 24'h4faf7e;
          13'h150C : pic_data = 24'h4faf82;
          13'h150D : pic_data = 24'h4faf89;
          13'h150E : pic_data = 24'h4faf8b;
          13'h150F : pic_data = 24'h4faf93;
          13'h1510 : pic_data = 24'h4faf9a;
          13'h1511 : pic_data = 24'h4faf9e;
          13'h1512 : pic_data = 24'h4fafa6;
          13'h1513 : pic_data = 24'h4fafa7;
          13'h1514 : pic_data = 24'h4fb0b0;
          13'h1515 : pic_data = 24'h4fa7af;
          13'h1516 : pic_data = 24'h4fa4af;
          13'h1517 : pic_data = 24'h4f9baf;
          13'h1518 : pic_data = 24'h4f95af;
          13'h1519 : pic_data = 24'h4f93af;
          13'h151A : pic_data = 24'h4f8caf;
          13'h151B : pic_data = 24'h4f87af;
          13'h151C : pic_data = 24'h4f80af;
          13'h151D : pic_data = 24'h4f78af;
          13'h151E : pic_data = 24'h4f76af;
          13'h151F : pic_data = 24'h4f6eaf;
          13'h1520 : pic_data = 24'h4f6aaf;
          13'h1521 : pic_data = 24'h4f63af;
          13'h1522 : pic_data = 24'h4f5baf;
          13'h1523 : pic_data = 24'h4f59af;
          13'h1524 : pic_data = 24'h4f52af;
          13'h1525 : pic_data = 24'h504faf;
          13'h1526 : pic_data = 24'h594faf;
          13'h1527 : pic_data = 24'h5f4faf;
          13'h1528 : pic_data = 24'h634faf;
          13'h1529 : pic_data = 24'h6c4faf;
          13'h152A : pic_data = 24'h6b4faf;
          13'h152B : pic_data = 24'h764faf;
          13'h152C : pic_data = 24'h7c4faf;
          13'h152D : pic_data = 24'h804faf;
          13'h152E : pic_data = 24'h8a4faf;
          13'h152F : pic_data = 24'h894faf;
          13'h1530 : pic_data = 24'h934faf;
          13'h1531 : pic_data = 24'h984faf;
          13'h1532 : pic_data = 24'h9c4faf;
          13'h1533 : pic_data = 24'ha64faf;
          13'h1534 : pic_data = 24'ha54faf;
          13'h1535 : pic_data = 24'hb04fb0;
          13'h1536 : pic_data = 24'haf4faa;
          13'h1537 : pic_data = 24'haf4fa5;
          13'h1538 : pic_data = 24'haf4f9b;
          13'h1539 : pic_data = 24'haf4f97;
          13'h153A : pic_data = 24'haf4f93;
          13'h153B : pic_data = 24'haf4f8e;
          13'h153C : pic_data = 24'haf4f89;
          13'h153D : pic_data = 24'haf4f7f;
          13'h153E : pic_data = 24'haf4f7a;
          13'h153F : pic_data = 24'haf4f75;
          13'h1540 : pic_data = 24'haf4f70;
          13'h1541 : pic_data = 24'haf4f6c;
          13'h1542 : pic_data = 24'haf4f62;
          13'h1543 : pic_data = 24'haf4f5e;
          13'h1544 : pic_data = 24'haf4f58;
          13'h1545 : pic_data = 24'had5051;
          13'h1546 : pic_data = 24'had5551;
          13'h1547 : pic_data = 24'had5951;
          13'h1548 : pic_data = 24'had6451;
          13'h1549 : pic_data = 24'had6851;
          13'h154A : pic_data = 24'had6b51;
          13'h154B : pic_data = 24'had7151;
          13'h154C : pic_data = 24'had7551;
          13'h154D : pic_data = 24'had8051;
          13'h154E : pic_data = 24'had8351;
          13'h154F : pic_data = 24'had8951;
          13'h1550 : pic_data = 24'had8c51;
          13'h1551 : pic_data = 24'had9251;
          13'h1552 : pic_data = 24'had9a51;
          13'h1553 : pic_data = 24'had9e51;
          13'h1554 : pic_data = 24'hada551;
          13'h1555 : pic_data = 24'hada851;
          13'h1556 : pic_data = 24'haeae51;
          13'h1557 : pic_data = 24'ha5ad51;
          13'h1558 : pic_data = 24'ha0ad51;
          13'h1559 : pic_data = 24'h9aad51;
          13'h155A : pic_data = 24'h93ad51;
          13'h155B : pic_data = 24'h93ad51;
          13'h155C : pic_data = 24'h89ad51;
          13'h155D : pic_data = 24'h86ad51;
          13'h155E : pic_data = 24'h80ad51;
          13'h155F : pic_data = 24'h76ad51;
          13'h1560 : pic_data = 24'h77ad51;
          13'h1561 : pic_data = 24'h6cad51;
          13'h1562 : pic_data = 24'h69ad51;
          13'h1563 : pic_data = 24'h64ad51;
          13'h1564 : pic_data = 24'h5bad51;
          13'h1565 : pic_data = 24'h5aad51;
          13'h1566 : pic_data = 24'h52ad50;
          13'h1567 : pic_data = 24'h50ad53;
          13'h1568 : pic_data = 24'h51ad59;
          13'h1569 : pic_data = 24'h51ad62;
          13'h156A : pic_data = 24'h51ad65;
          13'h156B : pic_data = 24'h51ad6c;
          13'h156C : pic_data = 24'h51ad6e;
          13'h156D : pic_data = 24'h51ad75;
          13'h156E : pic_data = 24'h51ad7e;
          13'h156F : pic_data = 24'h51ad82;
          13'h1570 : pic_data = 24'h51ad89;
          13'h1571 : pic_data = 24'h51ad8b;
          13'h1572 : pic_data = 24'h51ad93;
          13'h1573 : pic_data = 24'h51ad98;
          13'h1574 : pic_data = 24'h51ad9d;
          13'h1575 : pic_data = 24'h51ada5;
          13'h1576 : pic_data = 24'h51ada6;
          13'h1577 : pic_data = 24'h51aeae;
          13'h1578 : pic_data = 24'h51a6ad;
          13'h1579 : pic_data = 24'h51a3ad;
          13'h157A : pic_data = 24'h519aad;
          13'h157B : pic_data = 24'h5194ad;
          13'h157C : pic_data = 24'h5193ad;
          13'h157D : pic_data = 24'h518bad;
          13'h157E : pic_data = 24'h5187ad;
          13'h157F : pic_data = 24'h5180ad;
          13'h1580 : pic_data = 24'h5178ad;
          13'h1581 : pic_data = 24'h5176ad;
          13'h1582 : pic_data = 24'h516ead;
          13'h1583 : pic_data = 24'h516bad;
          13'h1584 : pic_data = 24'h5164ad;
          13'h1585 : pic_data = 24'h515cad;
          13'h1586 : pic_data = 24'h515aad;
          13'h1587 : pic_data = 24'h5153ad;
          13'h1588 : pic_data = 24'h5150ad;
          13'h1589 : pic_data = 24'h5a51ad;
          13'h158A : pic_data = 24'h6051ad;
          13'h158B : pic_data = 24'h6451ad;
          13'h158C : pic_data = 24'h6c51ad;
          13'h158D : pic_data = 24'h6c51ad;
          13'h158E : pic_data = 24'h7651ad;
          13'h158F : pic_data = 24'h7c51ad;
          13'h1590 : pic_data = 24'h8051ad;
          13'h1591 : pic_data = 24'h8951ad;
          13'h1592 : pic_data = 24'h8851ad;
          13'h1593 : pic_data = 24'h9351ad;
          13'h1594 : pic_data = 24'h9851ad;
          13'h1595 : pic_data = 24'h9b51ad;
          13'h1596 : pic_data = 24'ha551ad;
          13'h1597 : pic_data = 24'ha451ad;
          13'h1598 : pic_data = 24'hae51ae;
          13'h1599 : pic_data = 24'had51a8;
          13'h159A : pic_data = 24'had51a4;
          13'h159B : pic_data = 24'had519a;
          13'h159C : pic_data = 24'had5196;
          13'h159D : pic_data = 24'had5193;
          13'h159E : pic_data = 24'had518d;
          13'h159F : pic_data = 24'had5189;
          13'h15A0 : pic_data = 24'had517f;
          13'h15A1 : pic_data = 24'had517b;
          13'h15A2 : pic_data = 24'had5176;
          13'h15A3 : pic_data = 24'had5171;
          13'h15A4 : pic_data = 24'had516c;
          13'h15A5 : pic_data = 24'had5163;
          13'h15A6 : pic_data = 24'had515f;
          13'h15A7 : pic_data = 24'had5159;
          13'h15A8 : pic_data = 24'hae5050;
          13'h15A9 : pic_data = 24'hae5450;
          13'h15AA : pic_data = 24'hae5950;
          13'h15AB : pic_data = 24'hae6450;
          13'h15AC : pic_data = 24'hae6750;
          13'h15AD : pic_data = 24'hae6b50;
          13'h15AE : pic_data = 24'hae7050;
          13'h15AF : pic_data = 24'hae7550;
          13'h15B0 : pic_data = 24'hae8050;
          13'h15B1 : pic_data = 24'hae8350;
          13'h15B2 : pic_data = 24'hae8950;
          13'h15B3 : pic_data = 24'hae8c50;
          13'h15B4 : pic_data = 24'hae9350;
          13'h15B5 : pic_data = 24'hae9a50;
          13'h15B6 : pic_data = 24'hae9f50;
          13'h15B7 : pic_data = 24'haea550;
          13'h15B8 : pic_data = 24'haea950;
          13'h15B9 : pic_data = 24'hafae50;
          13'h15BA : pic_data = 24'ha5ae50;
          13'h15BB : pic_data = 24'ha1ae50;
          13'h15BC : pic_data = 24'h9bae50;
          13'h15BD : pic_data = 24'h93ae50;
          13'h15BE : pic_data = 24'h94ae50;
          13'h15BF : pic_data = 24'h89ae50;
          13'h15C0 : pic_data = 24'h86ae50;
          13'h15C1 : pic_data = 24'h80ae50;
          13'h15C2 : pic_data = 24'h75ae50;
          13'h15C3 : pic_data = 24'h76ae50;
          13'h15C4 : pic_data = 24'h6cae50;
          13'h15C5 : pic_data = 24'h68ae50;
          13'h15C6 : pic_data = 24'h64ae50;
          13'h15C7 : pic_data = 24'h5bae50;
          13'h15C8 : pic_data = 24'h5aae50;
          13'h15C9 : pic_data = 24'h52ae50;
          13'h15CA : pic_data = 24'h50ae53;
          13'h15CB : pic_data = 24'h50ae59;
          13'h15CC : pic_data = 24'h50ae62;
          13'h15CD : pic_data = 24'h50ae65;
          13'h15CE : pic_data = 24'h50ae6c;
          13'h15CF : pic_data = 24'h50ae6e;
          13'h15D0 : pic_data = 24'h50ae75;
          13'h15D1 : pic_data = 24'h50ae7e;
          13'h15D2 : pic_data = 24'h50ae82;
          13'h15D3 : pic_data = 24'h50ae89;
          13'h15D4 : pic_data = 24'h50ae8b;
          13'h15D5 : pic_data = 24'h50ae93;
          13'h15D6 : pic_data = 24'h50ae99;
          13'h15D7 : pic_data = 24'h50ae9d;
          13'h15D8 : pic_data = 24'h50aea5;
          13'h15D9 : pic_data = 24'h50aea6;
          13'h15DA : pic_data = 24'h50afaf;
          13'h15DB : pic_data = 24'h50a6ae;
          13'h15DC : pic_data = 24'h50a3ae;
          13'h15DD : pic_data = 24'h509aae;
          13'h15DE : pic_data = 24'h5094ae;
          13'h15DF : pic_data = 24'h5093ae;
          13'h15E0 : pic_data = 24'h508bae;
          13'h15E1 : pic_data = 24'h5087ae;
          13'h15E2 : pic_data = 24'h5080ae;
          13'h15E3 : pic_data = 24'h5078ae;
          13'h15E4 : pic_data = 24'h5076ae;
          13'h15E5 : pic_data = 24'h506eae;
          13'h15E6 : pic_data = 24'h506bae;
          13'h15E7 : pic_data = 24'h5063ae;
          13'h15E8 : pic_data = 24'h505cae;
          13'h15E9 : pic_data = 24'h505aae;
          13'h15EA : pic_data = 24'h5053ae;
          13'h15EB : pic_data = 24'h5050ae;
          13'h15EC : pic_data = 24'h5950ae;
          13'h15ED : pic_data = 24'h5f50ae;
          13'h15EE : pic_data = 24'h6450ae;
          13'h15EF : pic_data = 24'h6c50ae;
          13'h15F0 : pic_data = 24'h6b50ae;
          13'h15F1 : pic_data = 24'h7650ae;
          13'h15F2 : pic_data = 24'h7c50ae;
          13'h15F3 : pic_data = 24'h8050ae;
          13'h15F4 : pic_data = 24'h8950ae;
          13'h15F5 : pic_data = 24'h8950ae;
          13'h15F6 : pic_data = 24'h9350ae;
          13'h15F7 : pic_data = 24'h9850ae;
          13'h15F8 : pic_data = 24'h9b50ae;
          13'h15F9 : pic_data = 24'ha650ae;
          13'h15FA : pic_data = 24'ha550ae;
          13'h15FB : pic_data = 24'haf50ae;
          13'h15FC : pic_data = 24'hae50a9;
          13'h15FD : pic_data = 24'hae50a4;
          13'h15FE : pic_data = 24'hae509a;
          13'h15FF : pic_data = 24'hae5097;
          13'h1600 : pic_data = 24'hae5093;
          13'h1601 : pic_data = 24'hae508e;
          13'h1602 : pic_data = 24'hae5089;
          13'h1603 : pic_data = 24'hae507f;
          13'h1604 : pic_data = 24'hae507b;
          13'h1605 : pic_data = 24'hae5075;
          13'h1606 : pic_data = 24'hae5070;
          13'h1607 : pic_data = 24'hae506c;
          13'h1608 : pic_data = 24'hae5063;
          13'h1609 : pic_data = 24'hae505e;
          13'h160A : pic_data = 24'hae5059;
          13'h160B : pic_data = 24'hab5353;
          13'h160C : pic_data = 24'hab5753;
          13'h160D : pic_data = 24'hab5c53;
          13'h160E : pic_data = 24'hab6553;
          13'h160F : pic_data = 24'hab6953;
          13'h1610 : pic_data = 24'hab6e53;
          13'h1611 : pic_data = 24'hab7253;
          13'h1612 : pic_data = 24'hab7653;
          13'h1613 : pic_data = 24'hab8053;
          13'h1614 : pic_data = 24'hab8353;
          13'h1615 : pic_data = 24'hab8853;
          13'h1616 : pic_data = 24'hab8c53;
          13'h1617 : pic_data = 24'hab9153;
          13'h1618 : pic_data = 24'hab9853;
          13'h1619 : pic_data = 24'hab9d53;
          13'h161A : pic_data = 24'haba353;
          13'h161B : pic_data = 24'haba653;
          13'h161C : pic_data = 24'hacab53;
          13'h161D : pic_data = 24'ha3ab53;
          13'h161E : pic_data = 24'h9fab53;
          13'h161F : pic_data = 24'h99ab53;
          13'h1620 : pic_data = 24'h91ab53;
          13'h1621 : pic_data = 24'h92ab53;
          13'h1622 : pic_data = 24'h88ab53;
          13'h1623 : pic_data = 24'h85ab53;
          13'h1624 : pic_data = 24'h80ab53;
          13'h1625 : pic_data = 24'h76ab53;
          13'h1626 : pic_data = 24'h77ab53;
          13'h1627 : pic_data = 24'h6eab53;
          13'h1628 : pic_data = 24'h6bab53;
          13'h1629 : pic_data = 24'h65ab53;
          13'h162A : pic_data = 24'h5dab53;
          13'h162B : pic_data = 24'h5dab53;
          13'h162C : pic_data = 24'h55ab53;
          13'h162D : pic_data = 24'h53ab56;
          13'h162E : pic_data = 24'h53ab5c;
          13'h162F : pic_data = 24'h53ab64;
          13'h1630 : pic_data = 24'h53ab67;
          13'h1631 : pic_data = 24'h53ab6e;
          13'h1632 : pic_data = 24'h53ab6f;
          13'h1633 : pic_data = 24'h53ab76;
          13'h1634 : pic_data = 24'h53ab7e;
          13'h1635 : pic_data = 24'h53ab82;
          13'h1636 : pic_data = 24'h53ab88;
          13'h1637 : pic_data = 24'h53ab8a;
          13'h1638 : pic_data = 24'h53ab91;
          13'h1639 : pic_data = 24'h53ab97;
          13'h163A : pic_data = 24'h53ab9b;
          13'h163B : pic_data = 24'h53aba3;
          13'h163C : pic_data = 24'h53aba4;
          13'h163D : pic_data = 24'h53acac;
          13'h163E : pic_data = 24'h53a4ab;
          13'h163F : pic_data = 24'h53a1ab;
          13'h1640 : pic_data = 24'h5399ab;
          13'h1641 : pic_data = 24'h5393ab;
          13'h1642 : pic_data = 24'h5392ab;
          13'h1643 : pic_data = 24'h538bab;
          13'h1644 : pic_data = 24'h5386ab;
          13'h1645 : pic_data = 24'h5380ab;
          13'h1646 : pic_data = 24'h5379ab;
          13'h1647 : pic_data = 24'h5377ab;
          13'h1648 : pic_data = 24'h5370ab;
          13'h1649 : pic_data = 24'h536cab;
          13'h164A : pic_data = 24'h5365ab;
          13'h164B : pic_data = 24'h535fab;
          13'h164C : pic_data = 24'h535dab;
          13'h164D : pic_data = 24'h5356ab;
          13'h164E : pic_data = 24'h5353ab;
          13'h164F : pic_data = 24'h5d53ab;
          13'h1650 : pic_data = 24'h6253ab;
          13'h1651 : pic_data = 24'h6553ab;
          13'h1652 : pic_data = 24'h6e53ab;
          13'h1653 : pic_data = 24'h6e53ab;
          13'h1654 : pic_data = 24'h7653ab;
          13'h1655 : pic_data = 24'h7c53ab;
          13'h1656 : pic_data = 24'h8053ab;
          13'h1657 : pic_data = 24'h8953ab;
          13'h1658 : pic_data = 24'h8853ab;
          13'h1659 : pic_data = 24'h9253ab;
          13'h165A : pic_data = 24'h9653ab;
          13'h165B : pic_data = 24'h9a53ab;
          13'h165C : pic_data = 24'ha353ab;
          13'h165D : pic_data = 24'ha353ab;
          13'h165E : pic_data = 24'hac53ab;
          13'h165F : pic_data = 24'hab53a6;
          13'h1660 : pic_data = 24'hab53a2;
          13'h1661 : pic_data = 24'hab5399;
          13'h1662 : pic_data = 24'hab5395;
          13'h1663 : pic_data = 24'hab5391;
          13'h1664 : pic_data = 24'hab538c;
          13'h1665 : pic_data = 24'hab5388;
          13'h1666 : pic_data = 24'hab537f;
          13'h1667 : pic_data = 24'hab537a;
          13'h1668 : pic_data = 24'hab5376;
          13'h1669 : pic_data = 24'hab5372;
          13'h166A : pic_data = 24'hab536e;
          13'h166B : pic_data = 24'hab5364;
          13'h166C : pic_data = 24'hab5361;
          13'h166D : pic_data = 24'hab535c;
          13'h166E : pic_data = 24'ha95455;
          13'h166F : pic_data = 24'ha95955;
          13'h1670 : pic_data = 24'ha95d55;
          13'h1671 : pic_data = 24'ha96655;
          13'h1672 : pic_data = 24'ha96955;
          13'h1673 : pic_data = 24'ha96f55;
          13'h1674 : pic_data = 24'ha97355;
          13'h1675 : pic_data = 24'ha97655;
          13'h1676 : pic_data = 24'ha98055;
          13'h1677 : pic_data = 24'ha98455;
          13'h1678 : pic_data = 24'ha98755;
          13'h1679 : pic_data = 24'ha98b55;
          13'h167A : pic_data = 24'ha99055;
          13'h167B : pic_data = 24'ha99855;
          13'h167C : pic_data = 24'ha99c55;
          13'h167D : pic_data = 24'ha9a255;
          13'h167E : pic_data = 24'ha9a455;
          13'h167F : pic_data = 24'haaaa55;
          13'h1680 : pic_data = 24'ha2a955;
          13'h1681 : pic_data = 24'h9da955;
          13'h1682 : pic_data = 24'h99a955;
          13'h1683 : pic_data = 24'h91a955;
          13'h1684 : pic_data = 24'h91a955;
          13'h1685 : pic_data = 24'h88a955;
          13'h1686 : pic_data = 24'h85a955;
          13'h1687 : pic_data = 24'h80a955;
          13'h1688 : pic_data = 24'h77a955;
          13'h1689 : pic_data = 24'h77a955;
          13'h168A : pic_data = 24'h6fa955;
          13'h168B : pic_data = 24'h6ca955;
          13'h168C : pic_data = 24'h66a955;
          13'h168D : pic_data = 24'h5ea955;
          13'h168E : pic_data = 24'h5ea955;
          13'h168F : pic_data = 24'h56a954;
          13'h1690 : pic_data = 24'h54a957;
          13'h1691 : pic_data = 24'h55a95e;
          13'h1692 : pic_data = 24'h55a965;
          13'h1693 : pic_data = 24'h55a968;
          13'h1694 : pic_data = 24'h55a96f;
          13'h1695 : pic_data = 24'h55a970;
          13'h1696 : pic_data = 24'h55a976;
          13'h1697 : pic_data = 24'h55a97e;
          13'h1698 : pic_data = 24'h55a981;
          13'h1699 : pic_data = 24'h55a988;
          13'h169A : pic_data = 24'h55a989;
          13'h169B : pic_data = 24'h55a991;
          13'h169C : pic_data = 24'h55a997;
          13'h169D : pic_data = 24'h55a99a;
          13'h169E : pic_data = 24'h55a9a2;
          13'h169F : pic_data = 24'h55a9a3;
          13'h16A0 : pic_data = 24'h55aaaa;
          13'h16A1 : pic_data = 24'h55a3a9;
          13'h16A2 : pic_data = 24'h55a0a9;
          13'h16A3 : pic_data = 24'h5598a9;
          13'h16A4 : pic_data = 24'h5592a9;
          13'h16A5 : pic_data = 24'h5591a9;
          13'h16A6 : pic_data = 24'h558aa9;
          13'h16A7 : pic_data = 24'h5586a9;
          13'h16A8 : pic_data = 24'h5580a9;
          13'h16A9 : pic_data = 24'h5579a9;
          13'h16AA : pic_data = 24'h5577a9;
          13'h16AB : pic_data = 24'h5570a9;
          13'h16AC : pic_data = 24'h556da9;
          13'h16AD : pic_data = 24'h5565a9;
          13'h16AE : pic_data = 24'h5560a9;
          13'h16AF : pic_data = 24'h555ea9;
          13'h16B0 : pic_data = 24'h5557a9;
          13'h16B1 : pic_data = 24'h5554a9;
          13'h16B2 : pic_data = 24'h5e55a9;
          13'h16B3 : pic_data = 24'h6355a9;
          13'h16B4 : pic_data = 24'h6655a9;
          13'h16B5 : pic_data = 24'h7055a9;
          13'h16B6 : pic_data = 24'h6f55a9;
          13'h16B7 : pic_data = 24'h7755a9;
          13'h16B8 : pic_data = 24'h7d55a9;
          13'h16B9 : pic_data = 24'h8055a9;
          13'h16BA : pic_data = 24'h8855a9;
          13'h16BB : pic_data = 24'h8855a9;
          13'h16BC : pic_data = 24'h9155a9;
          13'h16BD : pic_data = 24'h9655a9;
          13'h16BE : pic_data = 24'h9955a9;
          13'h16BF : pic_data = 24'ha255a9;
          13'h16C0 : pic_data = 24'ha255a9;
          13'h16C1 : pic_data = 24'haa55aa;
          13'h16C2 : pic_data = 24'ha955a4;
          13'h16C3 : pic_data = 24'ha955a1;
          13'h16C4 : pic_data = 24'ha95598;
          13'h16C5 : pic_data = 24'ha95594;
          13'h16C6 : pic_data = 24'ha95591;
          13'h16C7 : pic_data = 24'ha9558b;
          13'h16C8 : pic_data = 24'ha95588;
          13'h16C9 : pic_data = 24'ha9557f;
          13'h16CA : pic_data = 24'ha9557a;
          13'h16CB : pic_data = 24'ha95577;
          13'h16CC : pic_data = 24'ha95573;
          13'h16CD : pic_data = 24'ha9556f;
          13'h16CE : pic_data = 24'ha95565;
          13'h16CF : pic_data = 24'ha95562;
          13'h16D0 : pic_data = 24'ha9555d;
          13'h16D1 : pic_data = 24'haa5454;
          13'h16D2 : pic_data = 24'haa5854;
          13'h16D3 : pic_data = 24'haa5d54;
          13'h16D4 : pic_data = 24'haa6654;
          13'h16D5 : pic_data = 24'haa6954;
          13'h16D6 : pic_data = 24'haa6e54;
          13'h16D7 : pic_data = 24'haa7254;
          13'h16D8 : pic_data = 24'haa7654;
          13'h16D9 : pic_data = 24'haa8054;
          13'h16DA : pic_data = 24'haa8454;
          13'h16DB : pic_data = 24'haa8854;
          13'h16DC : pic_data = 24'haa8c54;
          13'h16DD : pic_data = 24'haa9054;
          13'h16DE : pic_data = 24'haa9854;
          13'h16DF : pic_data = 24'haa9d54;
          13'h16E0 : pic_data = 24'haaa254;
          13'h16E1 : pic_data = 24'haaa554;
          13'h16E2 : pic_data = 24'habaa54;
          13'h16E3 : pic_data = 24'ha3aa54;
          13'h16E4 : pic_data = 24'h9eaa54;
          13'h16E5 : pic_data = 24'h99aa54;
          13'h16E6 : pic_data = 24'h91aa54;
          13'h16E7 : pic_data = 24'h92aa54;
          13'h16E8 : pic_data = 24'h88aa54;
          13'h16E9 : pic_data = 24'h85aa54;
          13'h16EA : pic_data = 24'h80aa54;
          13'h16EB : pic_data = 24'h77aa54;
          13'h16EC : pic_data = 24'h77aa54;
          13'h16ED : pic_data = 24'h6faa54;
          13'h16EE : pic_data = 24'h6caa54;
          13'h16EF : pic_data = 24'h65aa54;
          13'h16F0 : pic_data = 24'h5eaa54;
          13'h16F1 : pic_data = 24'h5eaa54;
          13'h16F2 : pic_data = 24'h56aa54;
          13'h16F3 : pic_data = 24'h54aa57;
          13'h16F4 : pic_data = 24'h54aa5d;
          13'h16F5 : pic_data = 24'h54aa65;
          13'h16F6 : pic_data = 24'h54aa68;
          13'h16F7 : pic_data = 24'h54aa6f;
          13'h16F8 : pic_data = 24'h54aa70;
          13'h16F9 : pic_data = 24'h54aa76;
          13'h16FA : pic_data = 24'h54aa7e;
          13'h16FB : pic_data = 24'h54aa81;
          13'h16FC : pic_data = 24'h54aa88;
          13'h16FD : pic_data = 24'h54aa89;
          13'h16FE : pic_data = 24'h54aa91;
          13'h16FF : pic_data = 24'h54aa97;
          13'h1700 : pic_data = 24'h54aa9a;
          13'h1701 : pic_data = 24'h54aaa2;
          13'h1702 : pic_data = 24'h54aaa3;
          13'h1703 : pic_data = 24'h54abab;
          13'h1704 : pic_data = 24'h54a4aa;
          13'h1705 : pic_data = 24'h54a0aa;
          13'h1706 : pic_data = 24'h5499aa;
          13'h1707 : pic_data = 24'h5492aa;
          13'h1708 : pic_data = 24'h5491aa;
          13'h1709 : pic_data = 24'h548baa;
          13'h170A : pic_data = 24'h5486aa;
          13'h170B : pic_data = 24'h5480aa;
          13'h170C : pic_data = 24'h5479aa;
          13'h170D : pic_data = 24'h5477aa;
          13'h170E : pic_data = 24'h5470aa;
          13'h170F : pic_data = 24'h546daa;
          13'h1710 : pic_data = 24'h5465aa;
          13'h1711 : pic_data = 24'h5460aa;
          13'h1712 : pic_data = 24'h545eaa;
          13'h1713 : pic_data = 24'h5457aa;
          13'h1714 : pic_data = 24'h5454aa;
          13'h1715 : pic_data = 24'h5e54aa;
          13'h1716 : pic_data = 24'h6254aa;
          13'h1717 : pic_data = 24'h6654aa;
          13'h1718 : pic_data = 24'h6f54aa;
          13'h1719 : pic_data = 24'h6f54aa;
          13'h171A : pic_data = 24'h7754aa;
          13'h171B : pic_data = 24'h7d54aa;
          13'h171C : pic_data = 24'h8054aa;
          13'h171D : pic_data = 24'h8854aa;
          13'h171E : pic_data = 24'h8854aa;
          13'h171F : pic_data = 24'h9154aa;
          13'h1720 : pic_data = 24'h9654aa;
          13'h1721 : pic_data = 24'h9954aa;
          13'h1722 : pic_data = 24'ha354aa;
          13'h1723 : pic_data = 24'ha254aa;
          13'h1724 : pic_data = 24'hab54aa;
          13'h1725 : pic_data = 24'haa54a5;
          13'h1726 : pic_data = 24'haa54a1;
          13'h1727 : pic_data = 24'haa5498;
          13'h1728 : pic_data = 24'haa5495;
          13'h1729 : pic_data = 24'haa5491;
          13'h172A : pic_data = 24'haa548c;
          13'h172B : pic_data = 24'haa5488;
          13'h172C : pic_data = 24'haa547f;
          13'h172D : pic_data = 24'haa547a;
          13'h172E : pic_data = 24'haa5476;
          13'h172F : pic_data = 24'haa5472;
          13'h1730 : pic_data = 24'haa546f;
          13'h1731 : pic_data = 24'haa5465;
          13'h1732 : pic_data = 24'haa5461;
          13'h1733 : pic_data = 24'haa545d;
          13'h1734 : pic_data = 24'ha75757;
          13'h1735 : pic_data = 24'ha75b57;
          13'h1736 : pic_data = 24'ha75f57;
          13'h1737 : pic_data = 24'ha76757;
          13'h1738 : pic_data = 24'ha76b57;
          13'h1739 : pic_data = 24'ha77057;
          13'h173A : pic_data = 24'ha77357;
          13'h173B : pic_data = 24'ha77757;
          13'h173C : pic_data = 24'ha78057;
          13'h173D : pic_data = 24'ha78357;
          13'h173E : pic_data = 24'ha78757;
          13'h173F : pic_data = 24'ha78a57;
          13'h1740 : pic_data = 24'ha78e57;
          13'h1741 : pic_data = 24'ha79757;
          13'h1742 : pic_data = 24'ha79b57;
          13'h1743 : pic_data = 24'ha79f57;
          13'h1744 : pic_data = 24'ha7a257;
          13'h1745 : pic_data = 24'ha8a857;
          13'h1746 : pic_data = 24'ha0a757;
          13'h1747 : pic_data = 24'h9ca757;
          13'h1748 : pic_data = 24'h98a757;
          13'h1749 : pic_data = 24'h8fa757;
          13'h174A : pic_data = 24'h8fa757;
          13'h174B : pic_data = 24'h88a757;
          13'h174C : pic_data = 24'h84a757;
          13'h174D : pic_data = 24'h80a757;
          13'h174E : pic_data = 24'h77a757;
          13'h174F : pic_data = 24'h78a757;
          13'h1750 : pic_data = 24'h71a757;
          13'h1751 : pic_data = 24'h6da757;
          13'h1752 : pic_data = 24'h67a757;
          13'h1753 : pic_data = 24'h60a757;
          13'h1754 : pic_data = 24'h60a757;
          13'h1755 : pic_data = 24'h58a757;
          13'h1756 : pic_data = 24'h57a75a;
          13'h1757 : pic_data = 24'h57a75f;
          13'h1758 : pic_data = 24'h57a766;
          13'h1759 : pic_data = 24'h57a76a;
          13'h175A : pic_data = 24'h57a770;
          13'h175B : pic_data = 24'h57a771;
          13'h175C : pic_data = 24'h57a777;
          13'h175D : pic_data = 24'h57a77e;
          13'h175E : pic_data = 24'h57a781;
          13'h175F : pic_data = 24'h57a787;
          13'h1760 : pic_data = 24'h57a788;
          13'h1761 : pic_data = 24'h57a78e;
          13'h1762 : pic_data = 24'h57a796;
          13'h1763 : pic_data = 24'h57a799;
          13'h1764 : pic_data = 24'h57a79f;
          13'h1765 : pic_data = 24'h57a7a0;
          13'h1766 : pic_data = 24'h57a8a8;
          13'h1767 : pic_data = 24'h57a1a7;
          13'h1768 : pic_data = 24'h579da7;
          13'h1769 : pic_data = 24'h5797a7;
          13'h176A : pic_data = 24'h5790a7;
          13'h176B : pic_data = 24'h578fa7;
          13'h176C : pic_data = 24'h5789a7;
          13'h176D : pic_data = 24'h5786a7;
          13'h176E : pic_data = 24'h5780a7;
          13'h176F : pic_data = 24'h5779a7;
          13'h1770 : pic_data = 24'h5778a7;
          13'h1771 : pic_data = 24'h5772a7;
          13'h1772 : pic_data = 24'h576ea7;
          13'h1773 : pic_data = 24'h5767a7;
          13'h1774 : pic_data = 24'h5761a7;
          13'h1775 : pic_data = 24'h5760a7;
          13'h1776 : pic_data = 24'h575aa7;
          13'h1777 : pic_data = 24'h5757a7;
          13'h1778 : pic_data = 24'h6057a7;
          13'h1779 : pic_data = 24'h6557a7;
          13'h177A : pic_data = 24'h6757a7;
          13'h177B : pic_data = 24'h7157a7;
          13'h177C : pic_data = 24'h7057a7;
          13'h177D : pic_data = 24'h7757a7;
          13'h177E : pic_data = 24'h7d57a7;
          13'h177F : pic_data = 24'h8057a7;
          13'h1780 : pic_data = 24'h8857a7;
          13'h1781 : pic_data = 24'h8757a7;
          13'h1782 : pic_data = 24'h8f57a7;
          13'h1783 : pic_data = 24'h9457a7;
          13'h1784 : pic_data = 24'h9857a7;
          13'h1785 : pic_data = 24'ha057a7;
          13'h1786 : pic_data = 24'h9f57a7;
          13'h1787 : pic_data = 24'ha857a8;
          13'h1788 : pic_data = 24'ha757a2;
          13'h1789 : pic_data = 24'ha7579f;
          13'h178A : pic_data = 24'ha75797;
          13'h178B : pic_data = 24'ha75792;
          13'h178C : pic_data = 24'ha7578f;
          13'h178D : pic_data = 24'ha7578a;
          13'h178E : pic_data = 24'ha75787;
          13'h178F : pic_data = 24'ha7577f;
          13'h1790 : pic_data = 24'ha7577b;
          13'h1791 : pic_data = 24'ha75777;
          13'h1792 : pic_data = 24'ha75773;
          13'h1793 : pic_data = 24'ha75771;
          13'h1794 : pic_data = 24'ha75766;
          13'h1795 : pic_data = 24'ha75763;
          13'h1796 : pic_data = 24'ha7575f;
          13'h1797 : pic_data = 24'ha55859;
          13'h1798 : pic_data = 24'ha55d59;
          13'h1799 : pic_data = 24'ha56059;
          13'h179A : pic_data = 24'ha56859;
          13'h179B : pic_data = 24'ha56b59;
          13'h179C : pic_data = 24'ha57159;
          13'h179D : pic_data = 24'ha57359;
          13'h179E : pic_data = 24'ha57759;
          13'h179F : pic_data = 24'ha58059;
          13'h17A0 : pic_data = 24'ha58259;
          13'h17A1 : pic_data = 24'ha58759;
          13'h17A2 : pic_data = 24'ha58959;
          13'h17A3 : pic_data = 24'ha58d59;
          13'h17A4 : pic_data = 24'ha59659;
          13'h17A5 : pic_data = 24'ha59959;
          13'h17A6 : pic_data = 24'ha59d59;
          13'h17A7 : pic_data = 24'ha5a059;
          13'h17A8 : pic_data = 24'ha6a659;
          13'h17A9 : pic_data = 24'h9ea559;
          13'h17AA : pic_data = 24'h9aa559;
          13'h17AB : pic_data = 24'h97a559;
          13'h17AC : pic_data = 24'h8da559;
          13'h17AD : pic_data = 24'h8ea559;
          13'h17AE : pic_data = 24'h87a559;
          13'h17AF : pic_data = 24'h83a559;
          13'h17B0 : pic_data = 24'h80a559;
          13'h17B1 : pic_data = 24'h78a559;
          13'h17B2 : pic_data = 24'h78a559;
          13'h17B3 : pic_data = 24'h71a559;
          13'h17B4 : pic_data = 24'h6ea559;
          13'h17B5 : pic_data = 24'h68a559;
          13'h17B6 : pic_data = 24'h61a559;
          13'h17B7 : pic_data = 24'h61a559;
          13'h17B8 : pic_data = 24'h59a558;
          13'h17B9 : pic_data = 24'h59a55b;
          13'h17BA : pic_data = 24'h59a561;
          13'h17BB : pic_data = 24'h59a567;
          13'h17BC : pic_data = 24'h59a56a;
          13'h17BD : pic_data = 24'h59a571;
          13'h17BE : pic_data = 24'h59a572;
          13'h17BF : pic_data = 24'h59a577;
          13'h17C0 : pic_data = 24'h59a57e;
          13'h17C1 : pic_data = 24'h59a581;
          13'h17C2 : pic_data = 24'h59a587;
          13'h17C3 : pic_data = 24'h59a588;
          13'h17C4 : pic_data = 24'h59a58d;
          13'h17C5 : pic_data = 24'h59a595;
          13'h17C6 : pic_data = 24'h59a598;
          13'h17C7 : pic_data = 24'h59a59e;
          13'h17C8 : pic_data = 24'h59a59f;
          13'h17C9 : pic_data = 24'h59a6a6;
          13'h17CA : pic_data = 24'h599fa5;
          13'h17CB : pic_data = 24'h599ba5;
          13'h17CC : pic_data = 24'h5997a5;
          13'h17CD : pic_data = 24'h598fa5;
          13'h17CE : pic_data = 24'h598ea5;
          13'h17CF : pic_data = 24'h5988a5;
          13'h17D0 : pic_data = 24'h5986a5;
          13'h17D1 : pic_data = 24'h5980a5;
          13'h17D2 : pic_data = 24'h5979a5;
          13'h17D3 : pic_data = 24'h5978a5;
          13'h17D4 : pic_data = 24'h5972a5;
          13'h17D5 : pic_data = 24'h596fa5;
          13'h17D6 : pic_data = 24'h5967a5;
          13'h17D7 : pic_data = 24'h5962a5;
          13'h17D8 : pic_data = 24'h5961a5;
          13'h17D9 : pic_data = 24'h595ba5;
          13'h17DA : pic_data = 24'h5958a5;
          13'h17DB : pic_data = 24'h6159a5;
          13'h17DC : pic_data = 24'h6659a5;
          13'h17DD : pic_data = 24'h6859a5;
          13'h17DE : pic_data = 24'h7159a5;
          13'h17DF : pic_data = 24'h7159a5;
          13'h17E0 : pic_data = 24'h7859a5;
          13'h17E1 : pic_data = 24'h7d59a5;
          13'h17E2 : pic_data = 24'h8059a5;
          13'h17E3 : pic_data = 24'h8759a5;
          13'h17E4 : pic_data = 24'h8759a5;
          13'h17E5 : pic_data = 24'h8d59a5;
          13'h17E6 : pic_data = 24'h9259a5;
          13'h17E7 : pic_data = 24'h9759a5;
          13'h17E8 : pic_data = 24'h9e59a5;
          13'h17E9 : pic_data = 24'h9e59a5;
          13'h17EA : pic_data = 24'ha659a6;
          13'h17EB : pic_data = 24'ha559a0;
          13'h17EC : pic_data = 24'ha5599e;
          13'h17ED : pic_data = 24'ha55996;
          13'h17EE : pic_data = 24'ha55991;
          13'h17EF : pic_data = 24'ha5598d;
          13'h17F0 : pic_data = 24'ha55989;
          13'h17F1 : pic_data = 24'ha55987;
          13'h17F2 : pic_data = 24'ha5597f;
          13'h17F3 : pic_data = 24'ha5597c;
          13'h17F4 : pic_data = 24'ha55978;
          13'h17F5 : pic_data = 24'ha55973;
          13'h17F6 : pic_data = 24'ha55971;
          13'h17F7 : pic_data = 24'ha55967;
          13'h17F8 : pic_data = 24'ha55963;
          13'h17F9 : pic_data = 24'ha55960;
          13'h17FA : pic_data = 24'ha65858;
          13'h17FB : pic_data = 24'ha65c58;
          13'h17FC : pic_data = 24'ha66058;
          13'h17FD : pic_data = 24'ha66858;
          13'h17FE : pic_data = 24'ha66b58;
          13'h17FF : pic_data = 24'ha67158;
          13'h1800 : pic_data = 24'ha67358;
          13'h1801 : pic_data = 24'ha67758;
          13'h1802 : pic_data = 24'ha68058;
          13'h1803 : pic_data = 24'ha68258;
          13'h1804 : pic_data = 24'ha68758;
          13'h1805 : pic_data = 24'ha68958;
          13'h1806 : pic_data = 24'ha68d58;
          13'h1807 : pic_data = 24'ha69658;
          13'h1808 : pic_data = 24'ha69a58;
          13'h1809 : pic_data = 24'ha69e58;
          13'h180A : pic_data = 24'ha6a058;
          13'h180B : pic_data = 24'ha7a658;
          13'h180C : pic_data = 24'h9ea658;
          13'h180D : pic_data = 24'h9ba658;
          13'h180E : pic_data = 24'h97a658;
          13'h180F : pic_data = 24'h8ea658;
          13'h1810 : pic_data = 24'h8ea658;
          13'h1811 : pic_data = 24'h87a658;
          13'h1812 : pic_data = 24'h84a658;
          13'h1813 : pic_data = 24'h80a658;
          13'h1814 : pic_data = 24'h78a658;
          13'h1815 : pic_data = 24'h78a658;
          13'h1816 : pic_data = 24'h71a658;
          13'h1817 : pic_data = 24'h6ea658;
          13'h1818 : pic_data = 24'h67a658;
          13'h1819 : pic_data = 24'h61a658;
          13'h181A : pic_data = 24'h61a658;
          13'h181B : pic_data = 24'h58a658;
          13'h181C : pic_data = 24'h58a65b;
          13'h181D : pic_data = 24'h58a660;
          13'h181E : pic_data = 24'h58a667;
          13'h181F : pic_data = 24'h58a66a;
          13'h1820 : pic_data = 24'h58a671;
          13'h1821 : pic_data = 24'h58a672;
          13'h1822 : pic_data = 24'h58a677;
          13'h1823 : pic_data = 24'h58a67e;
          13'h1824 : pic_data = 24'h58a681;
          13'h1825 : pic_data = 24'h58a687;
          13'h1826 : pic_data = 24'h58a688;
          13'h1827 : pic_data = 24'h58a68d;
          13'h1828 : pic_data = 24'h58a695;
          13'h1829 : pic_data = 24'h58a699;
          13'h182A : pic_data = 24'h58a69e;
          13'h182B : pic_data = 24'h58a69f;
          13'h182C : pic_data = 24'h58a7a7;
          13'h182D : pic_data = 24'h589fa6;
          13'h182E : pic_data = 24'h589ca6;
          13'h182F : pic_data = 24'h5897a6;
          13'h1830 : pic_data = 24'h588fa6;
          13'h1831 : pic_data = 24'h588ea6;
          13'h1832 : pic_data = 24'h5888a6;
          13'h1833 : pic_data = 24'h5886a6;
          13'h1834 : pic_data = 24'h5880a6;
          13'h1835 : pic_data = 24'h5879a6;
          13'h1836 : pic_data = 24'h5878a6;
          13'h1837 : pic_data = 24'h5872a6;
          13'h1838 : pic_data = 24'h586fa6;
          13'h1839 : pic_data = 24'h5867a6;
          13'h183A : pic_data = 24'h5862a6;
          13'h183B : pic_data = 24'h5861a6;
          13'h183C : pic_data = 24'h585ba6;
          13'h183D : pic_data = 24'h5858a6;
          13'h183E : pic_data = 24'h6158a6;
          13'h183F : pic_data = 24'h6658a6;
          13'h1840 : pic_data = 24'h6858a6;
          13'h1841 : pic_data = 24'h7158a6;
          13'h1842 : pic_data = 24'h7158a6;
          13'h1843 : pic_data = 24'h7858a6;
          13'h1844 : pic_data = 24'h7d58a6;
          13'h1845 : pic_data = 24'h8058a6;
          13'h1846 : pic_data = 24'h8758a6;
          13'h1847 : pic_data = 24'h8758a6;
          13'h1848 : pic_data = 24'h8e58a6;
          13'h1849 : pic_data = 24'h9358a6;
          13'h184A : pic_data = 24'h9858a6;
          13'h184B : pic_data = 24'h9e58a6;
          13'h184C : pic_data = 24'h9e58a6;
          13'h184D : pic_data = 24'ha758a6;
          13'h184E : pic_data = 24'ha658a0;
          13'h184F : pic_data = 24'ha6589e;
          13'h1850 : pic_data = 24'ha65896;
          13'h1851 : pic_data = 24'ha65892;
          13'h1852 : pic_data = 24'ha6588e;
          13'h1853 : pic_data = 24'ha65889;
          13'h1854 : pic_data = 24'ha65887;
          13'h1855 : pic_data = 24'ha6587f;
          13'h1856 : pic_data = 24'ha6587c;
          13'h1857 : pic_data = 24'ha65877;
          13'h1858 : pic_data = 24'ha65873;
          13'h1859 : pic_data = 24'ha65871;
          13'h185A : pic_data = 24'ha65867;
          13'h185B : pic_data = 24'ha65863;
          13'h185C : pic_data = 24'ha65860;
          13'h185D : pic_data = 24'ha35b5c;
          13'h185E : pic_data = 24'ha35f5c;
          13'h185F : pic_data = 24'ha3625c;
          13'h1860 : pic_data = 24'ha36a5c;
          13'h1861 : pic_data = 24'ha36d5c;
          13'h1862 : pic_data = 24'ha3715c;
          13'h1863 : pic_data = 24'ha3745c;
          13'h1864 : pic_data = 24'ha3785c;
          13'h1865 : pic_data = 24'ha3805c;
          13'h1866 : pic_data = 24'ha3825c;
          13'h1867 : pic_data = 24'ha3865c;
          13'h1868 : pic_data = 24'ha3895c;
          13'h1869 : pic_data = 24'ha38c5c;
          13'h186A : pic_data = 24'ha3955c;
          13'h186B : pic_data = 24'ha3985c;
          13'h186C : pic_data = 24'ha39c5c;
          13'h186D : pic_data = 24'ha39e5c;
          13'h186E : pic_data = 24'ha4a45c;
          13'h186F : pic_data = 24'h9ca35c;
          13'h1870 : pic_data = 24'h99a35c;
          13'h1871 : pic_data = 24'h95a35c;
          13'h1872 : pic_data = 24'h8da35c;
          13'h1873 : pic_data = 24'h8da35c;
          13'h1874 : pic_data = 24'h87a35c;
          13'h1875 : pic_data = 24'h84a35c;
          13'h1876 : pic_data = 24'h80a35c;
          13'h1877 : pic_data = 24'h78a35c;
          13'h1878 : pic_data = 24'h79a35c;
          13'h1879 : pic_data = 24'h72a35c;
          13'h187A : pic_data = 24'h6fa35c;
          13'h187B : pic_data = 24'h69a35c;
          13'h187C : pic_data = 24'h63a35c;
          13'h187D : pic_data = 24'h63a35c;
          13'h187E : pic_data = 24'h5ca35b;
          13'h187F : pic_data = 24'h5ca35e;
          13'h1880 : pic_data = 24'h5ca362;
          13'h1881 : pic_data = 24'h5ca369;
          13'h1882 : pic_data = 24'h5ca36c;
          13'h1883 : pic_data = 24'h5ca372;
          13'h1884 : pic_data = 24'h5ca373;
          13'h1885 : pic_data = 24'h5ca378;
          13'h1886 : pic_data = 24'h5ca37e;
          13'h1887 : pic_data = 24'h5ca381;
          13'h1888 : pic_data = 24'h5ca386;
          13'h1889 : pic_data = 24'h5ca387;
          13'h188A : pic_data = 24'h5ca38d;
          13'h188B : pic_data = 24'h5ca393;
          13'h188C : pic_data = 24'h5ca396;
          13'h188D : pic_data = 24'h5ca39c;
          13'h188E : pic_data = 24'h5ca39d;
          13'h188F : pic_data = 24'h5ca4a4;
          13'h1890 : pic_data = 24'h5c9da3;
          13'h1891 : pic_data = 24'h5c9aa3;
          13'h1892 : pic_data = 24'h5c95a3;
          13'h1893 : pic_data = 24'h5c8ea3;
          13'h1894 : pic_data = 24'h5c8da3;
          13'h1895 : pic_data = 24'h5c88a3;
          13'h1896 : pic_data = 24'h5c85a3;
          13'h1897 : pic_data = 24'h5c80a3;
          13'h1898 : pic_data = 24'h5c7aa3;
          13'h1899 : pic_data = 24'h5c79a3;
          13'h189A : pic_data = 24'h5c73a3;
          13'h189B : pic_data = 24'h5c70a3;
          13'h189C : pic_data = 24'h5c69a3;
          13'h189D : pic_data = 24'h5c64a3;
          13'h189E : pic_data = 24'h5c63a3;
          13'h189F : pic_data = 24'h5c5ea3;
          13'h18A0 : pic_data = 24'h5c5ba3;
          13'h18A1 : pic_data = 24'h625ca3;
          13'h18A2 : pic_data = 24'h685ca3;
          13'h18A3 : pic_data = 24'h6a5ca3;
          13'h18A4 : pic_data = 24'h725ca3;
          13'h18A5 : pic_data = 24'h725ca3;
          13'h18A6 : pic_data = 24'h785ca3;
          13'h18A7 : pic_data = 24'h7d5ca3;
          13'h18A8 : pic_data = 24'h805ca3;
          13'h18A9 : pic_data = 24'h865ca3;
          13'h18AA : pic_data = 24'h865ca3;
          13'h18AB : pic_data = 24'h8d5ca3;
          13'h18AC : pic_data = 24'h915ca3;
          13'h18AD : pic_data = 24'h955ca3;
          13'h18AE : pic_data = 24'h9c5ca3;
          13'h18AF : pic_data = 24'h9c5ca3;
          13'h18B0 : pic_data = 24'ha45ca4;
          13'h18B1 : pic_data = 24'ha35c9e;
          13'h18B2 : pic_data = 24'ha35c9c;
          13'h18B3 : pic_data = 24'ha35c94;
          13'h18B4 : pic_data = 24'ha35c90;
          13'h18B5 : pic_data = 24'ha35c8d;
          13'h18B6 : pic_data = 24'ha35c89;
          13'h18B7 : pic_data = 24'ha35c86;
          13'h18B8 : pic_data = 24'ha35c7f;
          13'h18B9 : pic_data = 24'ha35c7b;
          13'h18BA : pic_data = 24'ha35c78;
          13'h18BB : pic_data = 24'ha35c74;
          13'h18BC : pic_data = 24'ha35c72;
          13'h18BD : pic_data = 24'ha35c69;
          13'h18BE : pic_data = 24'ha35c65;
          13'h18BF : pic_data = 24'ha35c62;
          13'h18C0 : pic_data = 24'ha15d5e;
          13'h18C1 : pic_data = 24'ha1615e;
          13'h18C2 : pic_data = 24'ha1635e;
          13'h18C3 : pic_data = 24'ha16b5e;
          13'h18C4 : pic_data = 24'ha16d5e;
          13'h18C5 : pic_data = 24'ha1725e;
          13'h18C6 : pic_data = 24'ha1745e;
          13'h18C7 : pic_data = 24'ha1785e;
          13'h18C8 : pic_data = 24'ha1805e;
          13'h18C9 : pic_data = 24'ha1835e;
          13'h18CA : pic_data = 24'ha1855e;
          13'h18CB : pic_data = 24'ha1885e;
          13'h18CC : pic_data = 24'ha18c5e;
          13'h18CD : pic_data = 24'ha1945e;
          13'h18CE : pic_data = 24'ha1965e;
          13'h18CF : pic_data = 24'ha19b5e;
          13'h18D0 : pic_data = 24'ha19d5e;
          13'h18D1 : pic_data = 24'ha2a25e;
          13'h18D2 : pic_data = 24'h9ba15e;
          13'h18D3 : pic_data = 24'h97a15e;
          13'h18D4 : pic_data = 24'h94a15e;
          13'h18D5 : pic_data = 24'h8da15e;
          13'h18D6 : pic_data = 24'h8da15e;
          13'h18D7 : pic_data = 24'h86a15e;
          13'h18D8 : pic_data = 24'h84a15e;
          13'h18D9 : pic_data = 24'h80a15e;
          13'h18DA : pic_data = 24'h79a15e;
          13'h18DB : pic_data = 24'h79a15e;
          13'h18DC : pic_data = 24'h72a15e;
          13'h18DD : pic_data = 24'h70a15e;
          13'h18DE : pic_data = 24'h6ba15e;
          13'h18DF : pic_data = 24'h64a15e;
          13'h18E0 : pic_data = 24'h64a15e;
          13'h18E1 : pic_data = 24'h5ea15d;
          13'h18E2 : pic_data = 24'h5ea15f;
          13'h18E3 : pic_data = 24'h5ea163;
          13'h18E4 : pic_data = 24'h5ea16a;
          13'h18E5 : pic_data = 24'h5ea16c;
          13'h18E6 : pic_data = 24'h5ea172;
          13'h18E7 : pic_data = 24'h5ea173;
          13'h18E8 : pic_data = 24'h5ea178;
          13'h18E9 : pic_data = 24'h5ea17f;
          13'h18EA : pic_data = 24'h5ea181;
          13'h18EB : pic_data = 24'h5ea186;
          13'h18EC : pic_data = 24'h5ea187;
          13'h18ED : pic_data = 24'h5ea18c;
          13'h18EE : pic_data = 24'h5ea191;
          13'h18EF : pic_data = 24'h5ea195;
          13'h18F0 : pic_data = 24'h5ea19b;
          13'h18F1 : pic_data = 24'h5ea19c;
          13'h18F2 : pic_data = 24'h5ea2a2;
          13'h18F3 : pic_data = 24'h5e9ca1;
          13'h18F4 : pic_data = 24'h5e99a1;
          13'h18F5 : pic_data = 24'h5e93a1;
          13'h18F6 : pic_data = 24'h5e8ea1;
          13'h18F7 : pic_data = 24'h5e8da1;
          13'h18F8 : pic_data = 24'h5e87a1;
          13'h18F9 : pic_data = 24'h5e85a1;
          13'h18FA : pic_data = 24'h5e80a1;
          13'h18FB : pic_data = 24'h5e7aa1;
          13'h18FC : pic_data = 24'h5e79a1;
          13'h18FD : pic_data = 24'h5e73a1;
          13'h18FE : pic_data = 24'h5e71a1;
          13'h18FF : pic_data = 24'h5e6ba1;
          13'h1900 : pic_data = 24'h5e65a1;
          13'h1901 : pic_data = 24'h5e64a1;
          13'h1902 : pic_data = 24'h5e5fa1;
          13'h1903 : pic_data = 24'h5e5da1;
          13'h1904 : pic_data = 24'h645ea1;
          13'h1905 : pic_data = 24'h695ea1;
          13'h1906 : pic_data = 24'h6b5ea1;
          13'h1907 : pic_data = 24'h725ea1;
          13'h1908 : pic_data = 24'h725ea1;
          13'h1909 : pic_data = 24'h795ea1;
          13'h190A : pic_data = 24'h7d5ea1;
          13'h190B : pic_data = 24'h805ea1;
          13'h190C : pic_data = 24'h865ea1;
          13'h190D : pic_data = 24'h865ea1;
          13'h190E : pic_data = 24'h8d5ea1;
          13'h190F : pic_data = 24'h905ea1;
          13'h1910 : pic_data = 24'h945ea1;
          13'h1911 : pic_data = 24'h9b5ea1;
          13'h1912 : pic_data = 24'h9b5ea1;
          13'h1913 : pic_data = 24'ha25ea2;
          13'h1914 : pic_data = 24'ha15e9d;
          13'h1915 : pic_data = 24'ha15e9b;
          13'h1916 : pic_data = 24'ha15e93;
          13'h1917 : pic_data = 24'ha15e8f;
          13'h1918 : pic_data = 24'ha15e8d;
          13'h1919 : pic_data = 24'ha15e88;
          13'h191A : pic_data = 24'ha15e86;
          13'h191B : pic_data = 24'ha15e7f;
          13'h191C : pic_data = 24'ha15e7b;
          13'h191D : pic_data = 24'ha15e79;
          13'h191E : pic_data = 24'ha15e74;
          13'h191F : pic_data = 24'ha15e72;
          13'h1920 : pic_data = 24'ha15e6a;
          13'h1921 : pic_data = 24'ha15e66;
          13'h1922 : pic_data = 24'ha15e63;
          13'h1923 : pic_data = 24'ha25d5d;
          13'h1924 : pic_data = 24'ha2605d;
          13'h1925 : pic_data = 24'ha2635d;
          13'h1926 : pic_data = 24'ha26b5d;
          13'h1927 : pic_data = 24'ha26d5d;
          13'h1928 : pic_data = 24'ha2725d;
          13'h1929 : pic_data = 24'ha2745d;
          13'h192A : pic_data = 24'ha2785d;
          13'h192B : pic_data = 24'ha2805d;
          13'h192C : pic_data = 24'ha2835d;
          13'h192D : pic_data = 24'ha2865d;
          13'h192E : pic_data = 24'ha2885d;
          13'h192F : pic_data = 24'ha28c5d;
          13'h1930 : pic_data = 24'ha2945d;
          13'h1931 : pic_data = 24'ha2965d;
          13'h1932 : pic_data = 24'ha29b5d;
          13'h1933 : pic_data = 24'ha29d5d;
          13'h1934 : pic_data = 24'ha2a25d;
          13'h1935 : pic_data = 24'h9ba25d;
          13'h1936 : pic_data = 24'h98a25d;
          13'h1937 : pic_data = 24'h94a25d;
          13'h1938 : pic_data = 24'h8da25d;
          13'h1939 : pic_data = 24'h8da25d;
          13'h193A : pic_data = 24'h86a25d;
          13'h193B : pic_data = 24'h84a25d;
          13'h193C : pic_data = 24'h80a25d;
          13'h193D : pic_data = 24'h79a25d;
          13'h193E : pic_data = 24'h79a25d;
          13'h193F : pic_data = 24'h72a25d;
          13'h1940 : pic_data = 24'h70a25d;
          13'h1941 : pic_data = 24'h6ba25d;
          13'h1942 : pic_data = 24'h64a25d;
          13'h1943 : pic_data = 24'h64a25d;
          13'h1944 : pic_data = 24'h5ea25d;
          13'h1945 : pic_data = 24'h5da25f;
          13'h1946 : pic_data = 24'h5da263;
          13'h1947 : pic_data = 24'h5da26a;
          13'h1948 : pic_data = 24'h5da26c;
          13'h1949 : pic_data = 24'h5da272;
          13'h194A : pic_data = 24'h5da273;
          13'h194B : pic_data = 24'h5da278;
          13'h194C : pic_data = 24'h5da27f;
          13'h194D : pic_data = 24'h5da281;
          13'h194E : pic_data = 24'h5da286;
          13'h194F : pic_data = 24'h5da287;
          13'h1950 : pic_data = 24'h5da28d;
          13'h1951 : pic_data = 24'h5da292;
          13'h1952 : pic_data = 24'h5da295;
          13'h1953 : pic_data = 24'h5da29b;
          13'h1954 : pic_data = 24'h5da29c;
          13'h1955 : pic_data = 24'h5da2a2;
          13'h1956 : pic_data = 24'h5d9ca2;
          13'h1957 : pic_data = 24'h5d99a2;
          13'h1958 : pic_data = 24'h5d94a2;
          13'h1959 : pic_data = 24'h5d8ea2;
          13'h195A : pic_data = 24'h5d8da2;
          13'h195B : pic_data = 24'h5d87a2;
          13'h195C : pic_data = 24'h5d85a2;
          13'h195D : pic_data = 24'h5d80a2;
          13'h195E : pic_data = 24'h5d7aa2;
          13'h195F : pic_data = 24'h5d79a2;
          13'h1960 : pic_data = 24'h5d73a2;
          13'h1961 : pic_data = 24'h5d71a2;
          13'h1962 : pic_data = 24'h5d6aa2;
          13'h1963 : pic_data = 24'h5d65a2;
          13'h1964 : pic_data = 24'h5d64a2;
          13'h1965 : pic_data = 24'h5d5fa2;
          13'h1966 : pic_data = 24'h5e5da2;
          13'h1967 : pic_data = 24'h635da2;
          13'h1968 : pic_data = 24'h695da2;
          13'h1969 : pic_data = 24'h6b5da2;
          13'h196A : pic_data = 24'h725da2;
          13'h196B : pic_data = 24'h725da2;
          13'h196C : pic_data = 24'h795da2;
          13'h196D : pic_data = 24'h7d5da2;
          13'h196E : pic_data = 24'h805da2;
          13'h196F : pic_data = 24'h865da2;
          13'h1970 : pic_data = 24'h865da2;
          13'h1971 : pic_data = 24'h8d5da2;
          13'h1972 : pic_data = 24'h915da2;
          13'h1973 : pic_data = 24'h945da2;
          13'h1974 : pic_data = 24'h9b5da2;
          13'h1975 : pic_data = 24'h9b5da2;
          13'h1976 : pic_data = 24'ha25da2;
          13'h1977 : pic_data = 24'ha25d9d;
          13'h1978 : pic_data = 24'ha25d9b;
          13'h1979 : pic_data = 24'ha25d93;
          13'h197A : pic_data = 24'ha25d8f;
          13'h197B : pic_data = 24'ha25d8d;
          13'h197C : pic_data = 24'ha25d88;
          13'h197D : pic_data = 24'ha25d86;
          13'h197E : pic_data = 24'ha25d7f;
          13'h197F : pic_data = 24'ha25d7b;
          13'h1980 : pic_data = 24'ha25d79;
          13'h1981 : pic_data = 24'ha25d74;
          13'h1982 : pic_data = 24'ha25d72;
          13'h1983 : pic_data = 24'ha25d6a;
          13'h1984 : pic_data = 24'ha25d66;
          13'h1985 : pic_data = 24'ha25d63;
          13'h1986 : pic_data = 24'h9c6262;
          13'h1987 : pic_data = 24'h9c6562;
          13'h1988 : pic_data = 24'h9c6862;
          13'h1989 : pic_data = 24'h9c6d62;
          13'h198A : pic_data = 24'h9c7062;
          13'h198B : pic_data = 24'h9c7462;
          13'h198C : pic_data = 24'h9c7562;
          13'h198D : pic_data = 24'h9c7862;
          13'h198E : pic_data = 24'h9c8062;
          13'h198F : pic_data = 24'h9c8362;
          13'h1990 : pic_data = 24'h9c8662;
          13'h1991 : pic_data = 24'h9c8762;
          13'h1992 : pic_data = 24'h9c8a62;
          13'h1993 : pic_data = 24'h9c9262;
          13'h1994 : pic_data = 24'h9c9362;
          13'h1995 : pic_data = 24'h9c9662;
          13'h1996 : pic_data = 24'h9c9862;
          13'h1997 : pic_data = 24'h9d9c62;
          13'h1998 : pic_data = 24'h979c62;
          13'h1999 : pic_data = 24'h949c62;
          13'h199A : pic_data = 24'h929c62;
          13'h199B : pic_data = 24'h8b9c62;
          13'h199C : pic_data = 24'h8b9c62;
          13'h199D : pic_data = 24'h869c62;
          13'h199E : pic_data = 24'h849c62;
          13'h199F : pic_data = 24'h809c62;
          13'h19A0 : pic_data = 24'h799c62;
          13'h19A1 : pic_data = 24'h799c62;
          13'h19A2 : pic_data = 24'h759c62;
          13'h19A3 : pic_data = 24'h729c62;
          13'h19A4 : pic_data = 24'h6d9c62;
          13'h19A5 : pic_data = 24'h699c62;
          13'h19A6 : pic_data = 24'h689c62;
          13'h19A7 : pic_data = 24'h629c62;
          13'h19A8 : pic_data = 24'h629c64;
          13'h19A9 : pic_data = 24'h629c68;
          13'h19AA : pic_data = 24'h629c6c;
          13'h19AB : pic_data = 24'h629c6e;
          13'h19AC : pic_data = 24'h629c74;
          13'h19AD : pic_data = 24'h629c74;
          13'h19AE : pic_data = 24'h629c78;
          13'h19AF : pic_data = 24'h629c7f;
          13'h19B0 : pic_data = 24'h629c81;
          13'h19B1 : pic_data = 24'h629c86;
          13'h19B2 : pic_data = 24'h629c86;
          13'h19B3 : pic_data = 24'h629c8a;
          13'h19B4 : pic_data = 24'h629c90;
          13'h19B5 : pic_data = 24'h629c92;
          13'h19B6 : pic_data = 24'h629c96;
          13'h19B7 : pic_data = 24'h629c96;
          13'h19B8 : pic_data = 24'h629c9d;
          13'h19B9 : pic_data = 24'h62989c;
          13'h19BA : pic_data = 24'h62959c;
          13'h19BB : pic_data = 24'h62919c;
          13'h19BC : pic_data = 24'h628c9c;
          13'h19BD : pic_data = 24'h628b9c;
          13'h19BE : pic_data = 24'h62869c;
          13'h19BF : pic_data = 24'h62859c;
          13'h19C0 : pic_data = 24'h62809c;
          13'h19C1 : pic_data = 24'h627a9c;
          13'h19C2 : pic_data = 24'h62799c;
          13'h19C3 : pic_data = 24'h62769c;
          13'h19C4 : pic_data = 24'h62739c;
          13'h19C5 : pic_data = 24'h626c9c;
          13'h19C6 : pic_data = 24'h626a9c;
          13'h19C7 : pic_data = 24'h62689c;
          13'h19C8 : pic_data = 24'h62649c;
          13'h19C9 : pic_data = 24'h62629c;
          13'h19CA : pic_data = 24'h68629c;
          13'h19CB : pic_data = 24'h6b629c;
          13'h19CC : pic_data = 24'h6d629c;
          13'h19CD : pic_data = 24'h74629c;
          13'h19CE : pic_data = 24'h74629c;
          13'h19CF : pic_data = 24'h79629c;
          13'h19D0 : pic_data = 24'h7d629c;
          13'h19D1 : pic_data = 24'h80629c;
          13'h19D2 : pic_data = 24'h86629c;
          13'h19D3 : pic_data = 24'h86629c;
          13'h19D4 : pic_data = 24'h8a629c;
          13'h19D5 : pic_data = 24'h8e629c;
          13'h19D6 : pic_data = 24'h91629c;
          13'h19D7 : pic_data = 24'h97629c;
          13'h19D8 : pic_data = 24'h95629c;
          13'h19D9 : pic_data = 24'h9d629c;
          13'h19DA : pic_data = 24'h9c6299;
          13'h19DB : pic_data = 24'h9c6296;
          13'h19DC : pic_data = 24'h9c6291;
          13'h19DD : pic_data = 24'h9c628d;
          13'h19DE : pic_data = 24'h9c628a;
          13'h19DF : pic_data = 24'h9c6287;
          13'h19E0 : pic_data = 24'h9c6286;
          13'h19E1 : pic_data = 24'h9c627f;
          13'h19E2 : pic_data = 24'h9c627b;
          13'h19E3 : pic_data = 24'h9c6279;
          13'h19E4 : pic_data = 24'h9c6275;
          13'h19E5 : pic_data = 24'h9c6274;
          13'h19E6 : pic_data = 24'h9c626c;
          13'h19E7 : pic_data = 24'h9c626a;
          13'h19E8 : pic_data = 24'h9c6268;
          13'h19E9 : pic_data = 24'h9d6161;
          13'h19EA : pic_data = 24'h9d6461;
          13'h19EB : pic_data = 24'h9d6761;
          13'h19EC : pic_data = 24'h9d6d61;
          13'h19ED : pic_data = 24'h9d6f61;
          13'h19EE : pic_data = 24'h9d7461;
          13'h19EF : pic_data = 24'h9d7561;
          13'h19F0 : pic_data = 24'h9d7861;
          13'h19F1 : pic_data = 24'h9d8061;
          13'h19F2 : pic_data = 24'h9d8361;
          13'h19F3 : pic_data = 24'h9d8661;
          13'h19F4 : pic_data = 24'h9d8761;
          13'h19F5 : pic_data = 24'h9d8a61;
          13'h19F6 : pic_data = 24'h9d9261;
          13'h19F7 : pic_data = 24'h9d9361;
          13'h19F8 : pic_data = 24'h9d9761;
          13'h19F9 : pic_data = 24'h9d9861;
          13'h19FA : pic_data = 24'h9d9d61;
          13'h19FB : pic_data = 24'h979d61;
          13'h19FC : pic_data = 24'h959d61;
          13'h19FD : pic_data = 24'h929d61;
          13'h19FE : pic_data = 24'h8b9d61;
          13'h19FF : pic_data = 24'h8b9d61;
          13'h1A00 : pic_data = 24'h869d61;
          13'h1A01 : pic_data = 24'h849d61;
          13'h1A02 : pic_data = 24'h809d61;
          13'h1A03 : pic_data = 24'h799d61;
          13'h1A04 : pic_data = 24'h799d61;
          13'h1A05 : pic_data = 24'h749d61;
          13'h1A06 : pic_data = 24'h729d61;
          13'h1A07 : pic_data = 24'h6c9d61;
          13'h1A08 : pic_data = 24'h689d61;
          13'h1A09 : pic_data = 24'h689d61;
          13'h1A0A : pic_data = 24'h629d61;
          13'h1A0B : pic_data = 24'h619d63;
          13'h1A0C : pic_data = 24'h619d67;
          13'h1A0D : pic_data = 24'h619d6c;
          13'h1A0E : pic_data = 24'h619d6e;
          13'h1A0F : pic_data = 24'h619d74;
          13'h1A10 : pic_data = 24'h619d74;
          13'h1A11 : pic_data = 24'h619d78;
          13'h1A12 : pic_data = 24'h619d7f;
          13'h1A13 : pic_data = 24'h619d81;
          13'h1A14 : pic_data = 24'h619d86;
          13'h1A15 : pic_data = 24'h619d86;
          13'h1A16 : pic_data = 24'h619d8a;
          13'h1A17 : pic_data = 24'h619d90;
          13'h1A18 : pic_data = 24'h619d92;
          13'h1A19 : pic_data = 24'h619d97;
          13'h1A1A : pic_data = 24'h619d97;
          13'h1A1B : pic_data = 24'h619d9d;
          13'h1A1C : pic_data = 24'h61989d;
          13'h1A1D : pic_data = 24'h61969d;
          13'h1A1E : pic_data = 24'h61929d;
          13'h1A1F : pic_data = 24'h618c9d;
          13'h1A20 : pic_data = 24'h618b9d;
          13'h1A21 : pic_data = 24'h61869d;
          13'h1A22 : pic_data = 24'h61859d;
          13'h1A23 : pic_data = 24'h61809d;
          13'h1A24 : pic_data = 24'h617a9d;
          13'h1A25 : pic_data = 24'h61799d;
          13'h1A26 : pic_data = 24'h61759d;
          13'h1A27 : pic_data = 24'h61739d;
          13'h1A28 : pic_data = 24'h616c9d;
          13'h1A29 : pic_data = 24'h61699d;
          13'h1A2A : pic_data = 24'h61689d;
          13'h1A2B : pic_data = 24'h61639d;
          13'h1A2C : pic_data = 24'h62619d;
          13'h1A2D : pic_data = 24'h68619d;
          13'h1A2E : pic_data = 24'h6a619d;
          13'h1A2F : pic_data = 24'h6d619d;
          13'h1A30 : pic_data = 24'h74619d;
          13'h1A31 : pic_data = 24'h74619d;
          13'h1A32 : pic_data = 24'h78619d;
          13'h1A33 : pic_data = 24'h7c619d;
          13'h1A34 : pic_data = 24'h80619d;
          13'h1A35 : pic_data = 24'h86619d;
          13'h1A36 : pic_data = 24'h86619d;
          13'h1A37 : pic_data = 24'h8b619d;
          13'h1A38 : pic_data = 24'h8f619d;
          13'h1A39 : pic_data = 24'h91619d;
          13'h1A3A : pic_data = 24'h97619d;
          13'h1A3B : pic_data = 24'h96619d;
          13'h1A3C : pic_data = 24'h9d619d;
          13'h1A3D : pic_data = 24'h9d619a;
          13'h1A3E : pic_data = 24'h9d6197;
          13'h1A3F : pic_data = 24'h9d6191;
          13'h1A40 : pic_data = 24'h9d618d;
          13'h1A41 : pic_data = 24'h9d618b;
          13'h1A42 : pic_data = 24'h9d6187;
          13'h1A43 : pic_data = 24'h9d6186;
          13'h1A44 : pic_data = 24'h9d617f;
          13'h1A45 : pic_data = 24'h9d617b;
          13'h1A46 : pic_data = 24'h9d6178;
          13'h1A47 : pic_data = 24'h9d6175;
          13'h1A48 : pic_data = 24'h9d6174;
          13'h1A49 : pic_data = 24'h9d616c;
          13'h1A4A : pic_data = 24'h9d6169;
          13'h1A4B : pic_data = 24'h9d6167;
          13'h1A4C : pic_data = 24'h9d6161;
          13'h1A4D : pic_data = 24'h9d6461;
          13'h1A4E : pic_data = 24'h9d6761;
          13'h1A4F : pic_data = 24'h9d6d61;
          13'h1A50 : pic_data = 24'h9d6f61;
          13'h1A51 : pic_data = 24'h9d7461;
          13'h1A52 : pic_data = 24'h9d7561;
          13'h1A53 : pic_data = 24'h9d7861;
          13'h1A54 : pic_data = 24'h9d8061;
          13'h1A55 : pic_data = 24'h9d8361;
          13'h1A56 : pic_data = 24'h9d8661;
          13'h1A57 : pic_data = 24'h9d8761;
          13'h1A58 : pic_data = 24'h9d8a61;
          13'h1A59 : pic_data = 24'h9d9261;
          13'h1A5A : pic_data = 24'h9d9361;
          13'h1A5B : pic_data = 24'h9d9761;
          13'h1A5C : pic_data = 24'h9d9861;
          13'h1A5D : pic_data = 24'h9d9d61;
          13'h1A5E : pic_data = 24'h979d61;
          13'h1A5F : pic_data = 24'h959d61;
          13'h1A60 : pic_data = 24'h929d61;
          13'h1A61 : pic_data = 24'h8b9d61;
          13'h1A62 : pic_data = 24'h8b9d61;
          13'h1A63 : pic_data = 24'h869d61;
          13'h1A64 : pic_data = 24'h849d61;
          13'h1A65 : pic_data = 24'h809d61;
          13'h1A66 : pic_data = 24'h799d61;
          13'h1A67 : pic_data = 24'h799d61;
          13'h1A68 : pic_data = 24'h749d61;
          13'h1A69 : pic_data = 24'h729d61;
          13'h1A6A : pic_data = 24'h6c9d61;
          13'h1A6B : pic_data = 24'h689d61;
          13'h1A6C : pic_data = 24'h689d61;
          13'h1A6D : pic_data = 24'h629d61;
          13'h1A6E : pic_data = 24'h619d63;
          13'h1A6F : pic_data = 24'h619d67;
          13'h1A70 : pic_data = 24'h619d6b;
          13'h1A71 : pic_data = 24'h619d6e;
          13'h1A72 : pic_data = 24'h619d74;
          13'h1A73 : pic_data = 24'h619d74;
          13'h1A74 : pic_data = 24'h619d78;
          13'h1A75 : pic_data = 24'h619d7f;
          13'h1A76 : pic_data = 24'h619d81;
          13'h1A77 : pic_data = 24'h619d86;
          13'h1A78 : pic_data = 24'h619d86;
          13'h1A79 : pic_data = 24'h619d8a;
          13'h1A7A : pic_data = 24'h619d90;
          13'h1A7B : pic_data = 24'h619d92;
          13'h1A7C : pic_data = 24'h619d97;
          13'h1A7D : pic_data = 24'h619d97;
          13'h1A7E : pic_data = 24'h619d9d;
          13'h1A7F : pic_data = 24'h61999d;
          13'h1A80 : pic_data = 24'h61969d;
          13'h1A81 : pic_data = 24'h61929d;
          13'h1A82 : pic_data = 24'h618c9d;
          13'h1A83 : pic_data = 24'h618b9d;
          13'h1A84 : pic_data = 24'h61869d;
          13'h1A85 : pic_data = 24'h61859d;
          13'h1A86 : pic_data = 24'h61809d;
          13'h1A87 : pic_data = 24'h617a9d;
          13'h1A88 : pic_data = 24'h61799d;
          13'h1A89 : pic_data = 24'h61759d;
          13'h1A8A : pic_data = 24'h61739d;
          13'h1A8B : pic_data = 24'h616c9d;
          13'h1A8C : pic_data = 24'h61699d;
          13'h1A8D : pic_data = 24'h61689d;
          13'h1A8E : pic_data = 24'h61639d;
          13'h1A8F : pic_data = 24'h62619d;
          13'h1A90 : pic_data = 24'h68619d;
          13'h1A91 : pic_data = 24'h6a619d;
          13'h1A92 : pic_data = 24'h6d619d;
          13'h1A93 : pic_data = 24'h74619d;
          13'h1A94 : pic_data = 24'h74619d;
          13'h1A95 : pic_data = 24'h78619d;
          13'h1A96 : pic_data = 24'h7c619d;
          13'h1A97 : pic_data = 24'h80619d;
          13'h1A98 : pic_data = 24'h86619d;
          13'h1A99 : pic_data = 24'h86619d;
          13'h1A9A : pic_data = 24'h8b619d;
          13'h1A9B : pic_data = 24'h8f619d;
          13'h1A9C : pic_data = 24'h91619d;
          13'h1A9D : pic_data = 24'h97619d;
          13'h1A9E : pic_data = 24'h96619d;
          13'h1A9F : pic_data = 24'h9d619d;
          13'h1AA0 : pic_data = 24'h9d619a;
          13'h1AA1 : pic_data = 24'h9d6197;
          13'h1AA2 : pic_data = 24'h9d6192;
          13'h1AA3 : pic_data = 24'h9d618d;
          13'h1AA4 : pic_data = 24'h9d618b;
          13'h1AA5 : pic_data = 24'h9d6187;
          13'h1AA6 : pic_data = 24'h9d6186;
          13'h1AA7 : pic_data = 24'h9d617f;
          13'h1AA8 : pic_data = 24'h9d617b;
          13'h1AA9 : pic_data = 24'h9d6178;
          13'h1AAA : pic_data = 24'h9d6175;
          13'h1AAB : pic_data = 24'h9d6174;
          13'h1AAC : pic_data = 24'h9d616c;
          13'h1AAD : pic_data = 24'h9d6169;
          13'h1AAE : pic_data = 24'h9d6167;
          13'h1AAF : pic_data = 24'h986666;
          13'h1AB0 : pic_data = 24'h986866;
          13'h1AB1 : pic_data = 24'h986a66;
          13'h1AB2 : pic_data = 24'h987166;
          13'h1AB3 : pic_data = 24'h987366;
          13'h1AB4 : pic_data = 24'h987566;
          13'h1AB5 : pic_data = 24'h987666;
          13'h1AB6 : pic_data = 24'h987966;
          13'h1AB7 : pic_data = 24'h988066;
          13'h1AB8 : pic_data = 24'h988166;
          13'h1AB9 : pic_data = 24'h988566;
          13'h1ABA : pic_data = 24'h988666;
          13'h1ABB : pic_data = 24'h988966;
          13'h1ABC : pic_data = 24'h988d66;
          13'h1ABD : pic_data = 24'h989066;
          13'h1ABE : pic_data = 24'h989366;
          13'h1ABF : pic_data = 24'h989566;
          13'h1AC0 : pic_data = 24'h999866;
          13'h1AC1 : pic_data = 24'h939866;
          13'h1AC2 : pic_data = 24'h919866;
          13'h1AC3 : pic_data = 24'h8d9866;
          13'h1AC4 : pic_data = 24'h899866;
          13'h1AC5 : pic_data = 24'h8a9866;
          13'h1AC6 : pic_data = 24'h859866;
          13'h1AC7 : pic_data = 24'h829866;
          13'h1AC8 : pic_data = 24'h809866;
          13'h1AC9 : pic_data = 24'h7a9866;
          13'h1ACA : pic_data = 24'h7a9866;
          13'h1ACB : pic_data = 24'h759866;
          13'h1ACC : pic_data = 24'h749866;
          13'h1ACD : pic_data = 24'h719866;
          13'h1ACE : pic_data = 24'h6b9866;
          13'h1ACF : pic_data = 24'h6b9866;
          13'h1AD0 : pic_data = 24'h679866;
          13'h1AD1 : pic_data = 24'h669868;
          13'h1AD2 : pic_data = 24'h66986b;
          13'h1AD3 : pic_data = 24'h669870;
          13'h1AD4 : pic_data = 24'h669872;
          13'h1AD5 : pic_data = 24'h669875;
          13'h1AD6 : pic_data = 24'h669875;
          13'h1AD7 : pic_data = 24'h669879;
          13'h1AD8 : pic_data = 24'h66987f;
          13'h1AD9 : pic_data = 24'h669880;
          13'h1ADA : pic_data = 24'h669885;
          13'h1ADB : pic_data = 24'h669885;
          13'h1ADC : pic_data = 24'h66988a;
          13'h1ADD : pic_data = 24'h66988c;
          13'h1ADE : pic_data = 24'h66988f;
          13'h1ADF : pic_data = 24'h669894;
          13'h1AE0 : pic_data = 24'h669894;
          13'h1AE1 : pic_data = 24'h669999;
          13'h1AE2 : pic_data = 24'h669498;
          13'h1AE3 : pic_data = 24'h669398;
          13'h1AE4 : pic_data = 24'h668d98;
          13'h1AE5 : pic_data = 24'h668a98;
          13'h1AE6 : pic_data = 24'h668a98;
          13'h1AE7 : pic_data = 24'h668598;
          13'h1AE8 : pic_data = 24'h668498;
          13'h1AE9 : pic_data = 24'h668098;
          13'h1AEA : pic_data = 24'h667b98;
          13'h1AEB : pic_data = 24'h667a98;
          13'h1AEC : pic_data = 24'h667798;
          13'h1AED : pic_data = 24'h667498;
          13'h1AEE : pic_data = 24'h667198;
          13'h1AEF : pic_data = 24'h666d98;
          13'h1AF0 : pic_data = 24'h666b98;
          13'h1AF1 : pic_data = 24'h666898;
          13'h1AF2 : pic_data = 24'h676698;
          13'h1AF3 : pic_data = 24'h6b6698;
          13'h1AF4 : pic_data = 24'h6f6698;
          13'h1AF5 : pic_data = 24'h726698;
          13'h1AF6 : pic_data = 24'h756698;
          13'h1AF7 : pic_data = 24'h756698;
          13'h1AF8 : pic_data = 24'h7a6698;
          13'h1AF9 : pic_data = 24'h7e6698;
          13'h1AFA : pic_data = 24'h806698;
          13'h1AFB : pic_data = 24'h856698;
          13'h1AFC : pic_data = 24'h856698;
          13'h1AFD : pic_data = 24'h8a6698;
          13'h1AFE : pic_data = 24'h8b6698;
          13'h1AFF : pic_data = 24'h8e6698;
          13'h1B00 : pic_data = 24'h946698;
          13'h1B01 : pic_data = 24'h936698;
          13'h1B02 : pic_data = 24'h996698;
          13'h1B03 : pic_data = 24'h986695;
          13'h1B04 : pic_data = 24'h986694;
          13'h1B05 : pic_data = 24'h98668d;
          13'h1B06 : pic_data = 24'h98668b;
          13'h1B07 : pic_data = 24'h98668a;
          13'h1B08 : pic_data = 24'h986686;
          13'h1B09 : pic_data = 24'h986685;
          13'h1B0A : pic_data = 24'h98667f;
          13'h1B0B : pic_data = 24'h98667d;
          13'h1B0C : pic_data = 24'h98667a;
          13'h1B0D : pic_data = 24'h986676;
          13'h1B0E : pic_data = 24'h986675;
          13'h1B0F : pic_data = 24'h986671;
          13'h1B10 : pic_data = 24'h98666e;
          13'h1B11 : pic_data = 24'h98666a;
          13'h1B12 : pic_data = 24'h996565;
          13'h1B13 : pic_data = 24'h996765;
          13'h1B14 : pic_data = 24'h996a65;
          13'h1B15 : pic_data = 24'h997165;
          13'h1B16 : pic_data = 24'h997265;
          13'h1B17 : pic_data = 24'h997465;
          13'h1B18 : pic_data = 24'h997665;
          13'h1B19 : pic_data = 24'h997965;
          13'h1B1A : pic_data = 24'h998065;
          13'h1B1B : pic_data = 24'h998165;
          13'h1B1C : pic_data = 24'h998565;
          13'h1B1D : pic_data = 24'h998665;
          13'h1B1E : pic_data = 24'h998965;
          13'h1B1F : pic_data = 24'h998e65;
          13'h1B20 : pic_data = 24'h999165;
          13'h1B21 : pic_data = 24'h999465;
          13'h1B22 : pic_data = 24'h999565;
          13'h1B23 : pic_data = 24'h999965;
          13'h1B24 : pic_data = 24'h939965;
          13'h1B25 : pic_data = 24'h929965;
          13'h1B26 : pic_data = 24'h8e9965;
          13'h1B27 : pic_data = 24'h899965;
          13'h1B28 : pic_data = 24'h8a9965;
          13'h1B29 : pic_data = 24'h859965;
          13'h1B2A : pic_data = 24'h839965;
          13'h1B2B : pic_data = 24'h809965;
          13'h1B2C : pic_data = 24'h7a9965;
          13'h1B2D : pic_data = 24'h7a9965;
          13'h1B2E : pic_data = 24'h759965;
          13'h1B2F : pic_data = 24'h749965;
          13'h1B30 : pic_data = 24'h719965;
          13'h1B31 : pic_data = 24'h6b9965;
          13'h1B32 : pic_data = 24'h6b9965;
          13'h1B33 : pic_data = 24'h669965;
          13'h1B34 : pic_data = 24'h659967;
          13'h1B35 : pic_data = 24'h65996a;
          13'h1B36 : pic_data = 24'h659970;
          13'h1B37 : pic_data = 24'h659971;
          13'h1B38 : pic_data = 24'h659975;
          13'h1B39 : pic_data = 24'h659975;
          13'h1B3A : pic_data = 24'h659979;
          13'h1B3B : pic_data = 24'h65997f;
          13'h1B3C : pic_data = 24'h659980;
          13'h1B3D : pic_data = 24'h659985;
          13'h1B3E : pic_data = 24'h659985;
          13'h1B3F : pic_data = 24'h65998a;
          13'h1B40 : pic_data = 24'h65998d;
          13'h1B41 : pic_data = 24'h65998f;
          13'h1B42 : pic_data = 24'h659994;
          13'h1B43 : pic_data = 24'h659994;
          13'h1B44 : pic_data = 24'h659999;
          13'h1B45 : pic_data = 24'h659499;
          13'h1B46 : pic_data = 24'h659399;
          13'h1B47 : pic_data = 24'h658d99;
          13'h1B48 : pic_data = 24'h658a99;
          13'h1B49 : pic_data = 24'h658a99;
          13'h1B4A : pic_data = 24'h658599;
          13'h1B4B : pic_data = 24'h658499;
          13'h1B4C : pic_data = 24'h658099;
          13'h1B4D : pic_data = 24'h657b99;
          13'h1B4E : pic_data = 24'h657a99;
          13'h1B4F : pic_data = 24'h657699;
          13'h1B50 : pic_data = 24'h657399;
          13'h1B51 : pic_data = 24'h657199;
          13'h1B52 : pic_data = 24'h656c99;
          13'h1B53 : pic_data = 24'h656b99;
          13'h1B54 : pic_data = 24'h656799;
          13'h1B55 : pic_data = 24'h666599;
          13'h1B56 : pic_data = 24'h6a6599;
          13'h1B57 : pic_data = 24'h6f6599;
          13'h1B58 : pic_data = 24'h716599;
          13'h1B59 : pic_data = 24'h756599;
          13'h1B5A : pic_data = 24'h756599;
          13'h1B5B : pic_data = 24'h796599;
          13'h1B5C : pic_data = 24'h7e6599;
          13'h1B5D : pic_data = 24'h806599;
          13'h1B5E : pic_data = 24'h856599;
          13'h1B5F : pic_data = 24'h856599;
          13'h1B60 : pic_data = 24'h8a6599;
          13'h1B61 : pic_data = 24'h8b6599;
          13'h1B62 : pic_data = 24'h8e6599;
          13'h1B63 : pic_data = 24'h946599;
          13'h1B64 : pic_data = 24'h936599;
          13'h1B65 : pic_data = 24'h996599;
          13'h1B66 : pic_data = 24'h996595;
          13'h1B67 : pic_data = 24'h996594;
          13'h1B68 : pic_data = 24'h99658d;
          13'h1B69 : pic_data = 24'h99658c;
          13'h1B6A : pic_data = 24'h99658a;
          13'h1B6B : pic_data = 24'h996586;
          13'h1B6C : pic_data = 24'h996585;
          13'h1B6D : pic_data = 24'h99657f;
          13'h1B6E : pic_data = 24'h99657d;
          13'h1B6F : pic_data = 24'h996579;
          13'h1B70 : pic_data = 24'h996576;
          13'h1B71 : pic_data = 24'h996575;
          13'h1B72 : pic_data = 24'h996570;
          13'h1B73 : pic_data = 24'h99656d;
          13'h1B74 : pic_data = 24'h99656a;
          13'h1B75 : pic_data = 24'h996565;
          13'h1B76 : pic_data = 24'h996765;
          13'h1B77 : pic_data = 24'h996a65;
          13'h1B78 : pic_data = 24'h997165;
          13'h1B79 : pic_data = 24'h997265;
          13'h1B7A : pic_data = 24'h997465;
          13'h1B7B : pic_data = 24'h997665;
          13'h1B7C : pic_data = 24'h997965;
          13'h1B7D : pic_data = 24'h998065;
          13'h1B7E : pic_data = 24'h998165;
          13'h1B7F : pic_data = 24'h998565;
          13'h1B80 : pic_data = 24'h998665;
          13'h1B81 : pic_data = 24'h998965;
          13'h1B82 : pic_data = 24'h998e65;
          13'h1B83 : pic_data = 24'h999165;
          13'h1B84 : pic_data = 24'h999465;
          13'h1B85 : pic_data = 24'h999665;
          13'h1B86 : pic_data = 24'h999965;
          13'h1B87 : pic_data = 24'h939965;
          13'h1B88 : pic_data = 24'h929965;
          13'h1B89 : pic_data = 24'h8e9965;
          13'h1B8A : pic_data = 24'h899965;
          13'h1B8B : pic_data = 24'h8a9965;
          13'h1B8C : pic_data = 24'h859965;
          13'h1B8D : pic_data = 24'h839965;
          13'h1B8E : pic_data = 24'h809965;
          13'h1B8F : pic_data = 24'h7a9965;
          13'h1B90 : pic_data = 24'h7a9965;
          13'h1B91 : pic_data = 24'h759965;
          13'h1B92 : pic_data = 24'h749965;
          13'h1B93 : pic_data = 24'h719965;
          13'h1B94 : pic_data = 24'h6b9965;
          13'h1B95 : pic_data = 24'h6b9965;
          13'h1B96 : pic_data = 24'h669965;
          13'h1B97 : pic_data = 24'h659967;
          13'h1B98 : pic_data = 24'h65996a;
          13'h1B99 : pic_data = 24'h659970;
          13'h1B9A : pic_data = 24'h659971;
          13'h1B9B : pic_data = 24'h659975;
          13'h1B9C : pic_data = 24'h659975;
          13'h1B9D : pic_data = 24'h659979;
          13'h1B9E : pic_data = 24'h65997f;
          13'h1B9F : pic_data = 24'h659980;
          13'h1BA0 : pic_data = 24'h659985;
          13'h1BA1 : pic_data = 24'h659985;
          13'h1BA2 : pic_data = 24'h65998a;
          13'h1BA3 : pic_data = 24'h65998d;
          13'h1BA4 : pic_data = 24'h659990;
          13'h1BA5 : pic_data = 24'h659994;
          13'h1BA6 : pic_data = 24'h659994;
          13'h1BA7 : pic_data = 24'h659999;
          13'h1BA8 : pic_data = 24'h659499;
          13'h1BA9 : pic_data = 24'h659399;
          13'h1BAA : pic_data = 24'h658d99;
          13'h1BAB : pic_data = 24'h658a99;
          13'h1BAC : pic_data = 24'h658a99;
          13'h1BAD : pic_data = 24'h658599;
          13'h1BAE : pic_data = 24'h658499;
          13'h1BAF : pic_data = 24'h658099;
          13'h1BB0 : pic_data = 24'h657b99;
          13'h1BB1 : pic_data = 24'h657a99;
          13'h1BB2 : pic_data = 24'h657699;
          13'h1BB3 : pic_data = 24'h657399;
          13'h1BB4 : pic_data = 24'h657099;
          13'h1BB5 : pic_data = 24'h656c99;
          13'h1BB6 : pic_data = 24'h656a99;
          13'h1BB7 : pic_data = 24'h656799;
          13'h1BB8 : pic_data = 24'h666599;
          13'h1BB9 : pic_data = 24'h6a6599;
          13'h1BBA : pic_data = 24'h6e6599;
          13'h1BBB : pic_data = 24'h716599;
          13'h1BBC : pic_data = 24'h756599;
          13'h1BBD : pic_data = 24'h756599;
          13'h1BBE : pic_data = 24'h796599;
          13'h1BBF : pic_data = 24'h7e6599;
          13'h1BC0 : pic_data = 24'h806599;
          13'h1BC1 : pic_data = 24'h856599;
          13'h1BC2 : pic_data = 24'h856599;
          13'h1BC3 : pic_data = 24'h8a6599;
          13'h1BC4 : pic_data = 24'h8c6599;
          13'h1BC5 : pic_data = 24'h8e6599;
          13'h1BC6 : pic_data = 24'h946599;
          13'h1BC7 : pic_data = 24'h936599;
          13'h1BC8 : pic_data = 24'h996599;
          13'h1BC9 : pic_data = 24'h996596;
          13'h1BCA : pic_data = 24'h996594;
          13'h1BCB : pic_data = 24'h99658d;
          13'h1BCC : pic_data = 24'h99658c;
          13'h1BCD : pic_data = 24'h99658a;
          13'h1BCE : pic_data = 24'h996586;
          13'h1BCF : pic_data = 24'h996585;
          13'h1BD0 : pic_data = 24'h99657f;
          13'h1BD1 : pic_data = 24'h99657c;
          13'h1BD2 : pic_data = 24'h996579;
          13'h1BD3 : pic_data = 24'h996576;
          13'h1BD4 : pic_data = 24'h996575;
          13'h1BD5 : pic_data = 24'h996570;
          13'h1BD6 : pic_data = 24'h99656d;
          13'h1BD7 : pic_data = 24'h99656a;
          13'h1BD8 : pic_data = 24'h946a6a;
          13'h1BD9 : pic_data = 24'h946c6a;
          13'h1BDA : pic_data = 24'h946f6a;
          13'h1BDB : pic_data = 24'h94736a;
          13'h1BDC : pic_data = 24'h94756a;
          13'h1BDD : pic_data = 24'h94776a;
          13'h1BDE : pic_data = 24'h94796a;
          13'h1BDF : pic_data = 24'h947a6a;
          13'h1BE0 : pic_data = 24'h94806a;
          13'h1BE1 : pic_data = 24'h94826a;
          13'h1BE2 : pic_data = 24'h94836a;
          13'h1BE3 : pic_data = 24'h94856a;
          13'h1BE4 : pic_data = 24'h94876a;
          13'h1BE5 : pic_data = 24'h948c6a;
          13'h1BE6 : pic_data = 24'h948d6a;
          13'h1BE7 : pic_data = 24'h94906a;
          13'h1BE8 : pic_data = 24'h94926a;
          13'h1BE9 : pic_data = 24'h95946a;
          13'h1BEA : pic_data = 24'h90946a;
          13'h1BEB : pic_data = 24'h8e946a;
          13'h1BEC : pic_data = 24'h8b946a;
          13'h1BED : pic_data = 24'h87946a;
          13'h1BEE : pic_data = 24'h88946a;
          13'h1BEF : pic_data = 24'h83946a;
          13'h1BF0 : pic_data = 24'h81946a;
          13'h1BF1 : pic_data = 24'h80946a;
          13'h1BF2 : pic_data = 24'h7b946a;
          13'h1BF3 : pic_data = 24'h7b946a;
          13'h1BF4 : pic_data = 24'h78946a;
          13'h1BF5 : pic_data = 24'h76946a;
          13'h1BF6 : pic_data = 24'h73946a;
          13'h1BF7 : pic_data = 24'h70946a;
          13'h1BF8 : pic_data = 24'h6f946a;
          13'h1BF9 : pic_data = 24'h6b946a;
          13'h1BFA : pic_data = 24'h6a946c;
          13'h1BFB : pic_data = 24'h6a946f;
          13'h1BFC : pic_data = 24'h6a9472;
          13'h1BFD : pic_data = 24'h6a9474;
          13'h1BFE : pic_data = 24'h6a9477;
          13'h1BFF : pic_data = 24'h6a9477;
          13'h1C00 : pic_data = 24'h6a947a;
          13'h1C01 : pic_data = 24'h6a947f;
          13'h1C02 : pic_data = 24'h6a9480;
          13'h1C03 : pic_data = 24'h6a9484;
          13'h1C04 : pic_data = 24'h6a9484;
          13'h1C05 : pic_data = 24'h6a9487;
          13'h1C06 : pic_data = 24'h6a948a;
          13'h1C07 : pic_data = 24'h6a948c;
          13'h1C08 : pic_data = 24'h6a9491;
          13'h1C09 : pic_data = 24'h6a9491;
          13'h1C0A : pic_data = 24'h6a9494;
          13'h1C0B : pic_data = 24'h6a9194;
          13'h1C0C : pic_data = 24'h6a8f94;
          13'h1C0D : pic_data = 24'h6a8b94;
          13'h1C0E : pic_data = 24'h6a8894;
          13'h1C0F : pic_data = 24'h6a8894;
          13'h1C10 : pic_data = 24'h6a8494;
          13'h1C11 : pic_data = 24'h6a8394;
          13'h1C12 : pic_data = 24'h6a8094;
          13'h1C13 : pic_data = 24'h6a7b94;
          13'h1C14 : pic_data = 24'h6a7b94;
          13'h1C15 : pic_data = 24'h6a7794;
          13'h1C16 : pic_data = 24'h6a7694;
          13'h1C17 : pic_data = 24'h6a7394;
          13'h1C18 : pic_data = 24'h6a7094;
          13'h1C19 : pic_data = 24'h6a6f94;
          13'h1C1A : pic_data = 24'h6a6c94;
          13'h1C1B : pic_data = 24'h6b6a94;
          13'h1C1C : pic_data = 24'h6f6a94;
          13'h1C1D : pic_data = 24'h726a94;
          13'h1C1E : pic_data = 24'h746a94;
          13'h1C1F : pic_data = 24'h776a94;
          13'h1C20 : pic_data = 24'h776a94;
          13'h1C21 : pic_data = 24'h7b6a94;
          13'h1C22 : pic_data = 24'h7e6a94;
          13'h1C23 : pic_data = 24'h7f6a94;
          13'h1C24 : pic_data = 24'h846a94;
          13'h1C25 : pic_data = 24'h836a94;
          13'h1C26 : pic_data = 24'h886a94;
          13'h1C27 : pic_data = 24'h896a94;
          13'h1C28 : pic_data = 24'h8b6a94;
          13'h1C29 : pic_data = 24'h916a94;
          13'h1C2A : pic_data = 24'h906a94;
          13'h1C2B : pic_data = 24'h956a94;
          13'h1C2C : pic_data = 24'h946a92;
          13'h1C2D : pic_data = 24'h946a91;
          13'h1C2E : pic_data = 24'h946a8b;
          13'h1C2F : pic_data = 24'h946a89;
          13'h1C30 : pic_data = 24'h946a87;
          13'h1C31 : pic_data = 24'h946a85;
          13'h1C32 : pic_data = 24'h946a84;
          13'h1C33 : pic_data = 24'h946a7f;
          13'h1C34 : pic_data = 24'h946a7c;
          13'h1C35 : pic_data = 24'h946a7b;
          13'h1C36 : pic_data = 24'h946a79;
          13'h1C37 : pic_data = 24'h946a77;
          13'h1C38 : pic_data = 24'h946a72;
          13'h1C39 : pic_data = 24'h946a71;
          13'h1C3A : pic_data = 24'h946a6f;
          13'h1C3B : pic_data = 24'h956969;
          13'h1C3C : pic_data = 24'h956b69;
          13'h1C3D : pic_data = 24'h956e69;
          13'h1C3E : pic_data = 24'h957369;
          13'h1C3F : pic_data = 24'h957469;
          13'h1C40 : pic_data = 24'h957669;
          13'h1C41 : pic_data = 24'h957869;
          13'h1C42 : pic_data = 24'h957a69;
          13'h1C43 : pic_data = 24'h958069;
          13'h1C44 : pic_data = 24'h958269;
          13'h1C45 : pic_data = 24'h958469;
          13'h1C46 : pic_data = 24'h958669;
          13'h1C47 : pic_data = 24'h958769;
          13'h1C48 : pic_data = 24'h958c69;
          13'h1C49 : pic_data = 24'h958d69;
          13'h1C4A : pic_data = 24'h959169;
          13'h1C4B : pic_data = 24'h959369;
          13'h1C4C : pic_data = 24'h959569;
          13'h1C4D : pic_data = 24'h909569;
          13'h1C4E : pic_data = 24'h8f9569;
          13'h1C4F : pic_data = 24'h8c9569;
          13'h1C50 : pic_data = 24'h879569;
          13'h1C51 : pic_data = 24'h889569;
          13'h1C52 : pic_data = 24'h839569;
          13'h1C53 : pic_data = 24'h829569;
          13'h1C54 : pic_data = 24'h809569;
          13'h1C55 : pic_data = 24'h7b9569;
          13'h1C56 : pic_data = 24'h7b9569;
          13'h1C57 : pic_data = 24'h779569;
          13'h1C58 : pic_data = 24'h769569;
          13'h1C59 : pic_data = 24'h729569;
          13'h1C5A : pic_data = 24'h6f9569;
          13'h1C5B : pic_data = 24'h6f9569;
          13'h1C5C : pic_data = 24'h6a9569;
          13'h1C5D : pic_data = 24'h69956b;
          13'h1C5E : pic_data = 24'h69956e;
          13'h1C5F : pic_data = 24'h699572;
          13'h1C60 : pic_data = 24'h699573;
          13'h1C61 : pic_data = 24'h699577;
          13'h1C62 : pic_data = 24'h699577;
          13'h1C63 : pic_data = 24'h69957a;
          13'h1C64 : pic_data = 24'h69957f;
          13'h1C65 : pic_data = 24'h699580;
          13'h1C66 : pic_data = 24'h699584;
          13'h1C67 : pic_data = 24'h699584;
          13'h1C68 : pic_data = 24'h699588;
          13'h1C69 : pic_data = 24'h69958b;
          13'h1C6A : pic_data = 24'h69958c;
          13'h1C6B : pic_data = 24'h699591;
          13'h1C6C : pic_data = 24'h699591;
          13'h1C6D : pic_data = 24'h699595;
          13'h1C6E : pic_data = 24'h699195;
          13'h1C6F : pic_data = 24'h699095;
          13'h1C70 : pic_data = 24'h698b95;
          13'h1C71 : pic_data = 24'h698895;
          13'h1C72 : pic_data = 24'h698895;
          13'h1C73 : pic_data = 24'h698495;
          13'h1C74 : pic_data = 24'h698395;
          13'h1C75 : pic_data = 24'h698095;
          13'h1C76 : pic_data = 24'h697b95;
          13'h1C77 : pic_data = 24'h697b95;
          13'h1C78 : pic_data = 24'h697795;
          13'h1C79 : pic_data = 24'h697695;
          13'h1C7A : pic_data = 24'h697295;
          13'h1C7B : pic_data = 24'h696f95;
          13'h1C7C : pic_data = 24'h696f95;
          13'h1C7D : pic_data = 24'h696b95;
          13'h1C7E : pic_data = 24'h6a6995;
          13'h1C7F : pic_data = 24'h6f6995;
          13'h1C80 : pic_data = 24'h726995;
          13'h1C81 : pic_data = 24'h736995;
          13'h1C82 : pic_data = 24'h776995;
          13'h1C83 : pic_data = 24'h776995;
          13'h1C84 : pic_data = 24'h7a6995;
          13'h1C85 : pic_data = 24'h7e6995;
          13'h1C86 : pic_data = 24'h7f6995;
          13'h1C87 : pic_data = 24'h846995;
          13'h1C88 : pic_data = 24'h836995;
          13'h1C89 : pic_data = 24'h886995;
          13'h1C8A : pic_data = 24'h8a6995;
          13'h1C8B : pic_data = 24'h8b6995;
          13'h1C8C : pic_data = 24'h916995;
          13'h1C8D : pic_data = 24'h906995;
          13'h1C8E : pic_data = 24'h956995;
          13'h1C8F : pic_data = 24'h956993;
          13'h1C90 : pic_data = 24'h956991;
          13'h1C91 : pic_data = 24'h95698b;
          13'h1C92 : pic_data = 24'h95698a;
          13'h1C93 : pic_data = 24'h956988;
          13'h1C94 : pic_data = 24'h956986;
          13'h1C95 : pic_data = 24'h956984;
          13'h1C96 : pic_data = 24'h95697f;
          13'h1C97 : pic_data = 24'h95697c;
          13'h1C98 : pic_data = 24'h95697a;
          13'h1C99 : pic_data = 24'h956978;
          13'h1C9A : pic_data = 24'h956977;
          13'h1C9B : pic_data = 24'h956972;
          13'h1C9C : pic_data = 24'h956970;
          13'h1C9D : pic_data = 24'h95696e;
          13'h1C9E : pic_data = 24'h956969;
          13'h1C9F : pic_data = 24'h956b69;
          13'h1CA0 : pic_data = 24'h956e69;
          13'h1CA1 : pic_data = 24'h957369;
          13'h1CA2 : pic_data = 24'h957469;
          13'h1CA3 : pic_data = 24'h957669;
          13'h1CA4 : pic_data = 24'h957869;
          13'h1CA5 : pic_data = 24'h957a69;
          13'h1CA6 : pic_data = 24'h958069;
          13'h1CA7 : pic_data = 24'h958269;
          13'h1CA8 : pic_data = 24'h958469;
          13'h1CA9 : pic_data = 24'h958669;
          13'h1CAA : pic_data = 24'h958769;
          13'h1CAB : pic_data = 24'h958c69;
          13'h1CAC : pic_data = 24'h958e69;
          13'h1CAD : pic_data = 24'h959169;
          13'h1CAE : pic_data = 24'h959369;
          13'h1CAF : pic_data = 24'h959569;
          13'h1CB0 : pic_data = 24'h919569;
          13'h1CB1 : pic_data = 24'h8f9569;
          13'h1CB2 : pic_data = 24'h8c9569;
          13'h1CB3 : pic_data = 24'h879569;
          13'h1CB4 : pic_data = 24'h889569;
          13'h1CB5 : pic_data = 24'h839569;
          13'h1CB6 : pic_data = 24'h829569;
          13'h1CB7 : pic_data = 24'h809569;
          13'h1CB8 : pic_data = 24'h7b9569;
          13'h1CB9 : pic_data = 24'h7b9569;
          13'h1CBA : pic_data = 24'h779569;
          13'h1CBB : pic_data = 24'h759569;
          13'h1CBC : pic_data = 24'h729569;
          13'h1CBD : pic_data = 24'h6f9569;
          13'h1CBE : pic_data = 24'h6f9569;
          13'h1CBF : pic_data = 24'h6a9569;
          13'h1CC0 : pic_data = 24'h69956b;
          13'h1CC1 : pic_data = 24'h69956e;
          13'h1CC2 : pic_data = 24'h699571;
          13'h1CC3 : pic_data = 24'h699573;
          13'h1CC4 : pic_data = 24'h699577;
          13'h1CC5 : pic_data = 24'h699577;
          13'h1CC6 : pic_data = 24'h69957a;
          13'h1CC7 : pic_data = 24'h69957f;
          13'h1CC8 : pic_data = 24'h699580;
          13'h1CC9 : pic_data = 24'h699584;
          13'h1CCA : pic_data = 24'h699584;
          13'h1CCB : pic_data = 24'h699588;
          13'h1CCC : pic_data = 24'h69958b;
          13'h1CCD : pic_data = 24'h69958c;
          13'h1CCE : pic_data = 24'h699591;
          13'h1CCF : pic_data = 24'h699592;
          13'h1CD0 : pic_data = 24'h699595;
          13'h1CD1 : pic_data = 24'h699295;
          13'h1CD2 : pic_data = 24'h699095;
          13'h1CD3 : pic_data = 24'h698c95;
          13'h1CD4 : pic_data = 24'h698895;
          13'h1CD5 : pic_data = 24'h698895;
          13'h1CD6 : pic_data = 24'h698495;
          13'h1CD7 : pic_data = 24'h698395;
          13'h1CD8 : pic_data = 24'h698095;
          13'h1CD9 : pic_data = 24'h697b95;
          13'h1CDA : pic_data = 24'h697b95;
          13'h1CDB : pic_data = 24'h697795;
          13'h1CDC : pic_data = 24'h697595;
          13'h1CDD : pic_data = 24'h697295;
          13'h1CDE : pic_data = 24'h696f95;
          13'h1CDF : pic_data = 24'h696e95;
          13'h1CE0 : pic_data = 24'h696b95;
          13'h1CE1 : pic_data = 24'h6a6995;
          13'h1CE2 : pic_data = 24'h6e6995;
          13'h1CE3 : pic_data = 24'h716995;
          13'h1CE4 : pic_data = 24'h736995;
          13'h1CE5 : pic_data = 24'h776995;
          13'h1CE6 : pic_data = 24'h776995;
          13'h1CE7 : pic_data = 24'h7a6995;
          13'h1CE8 : pic_data = 24'h7e6995;
          13'h1CE9 : pic_data = 24'h7f6995;
          13'h1CEA : pic_data = 24'h846995;
          13'h1CEB : pic_data = 24'h836995;
          13'h1CEC : pic_data = 24'h886995;
          13'h1CED : pic_data = 24'h8a6995;
          13'h1CEE : pic_data = 24'h8b6995;
          13'h1CEF : pic_data = 24'h916995;
          13'h1CF0 : pic_data = 24'h906995;
          13'h1CF1 : pic_data = 24'h956995;
          13'h1CF2 : pic_data = 24'h956993;
          13'h1CF3 : pic_data = 24'h956991;
          13'h1CF4 : pic_data = 24'h95698b;
          13'h1CF5 : pic_data = 24'h95698a;
          13'h1CF6 : pic_data = 24'h956988;
          13'h1CF7 : pic_data = 24'h956986;
          13'h1CF8 : pic_data = 24'h956984;
          13'h1CF9 : pic_data = 24'h95697f;
          13'h1CFA : pic_data = 24'h95697c;
          13'h1CFB : pic_data = 24'h95697a;
          13'h1CFC : pic_data = 24'h956978;
          13'h1CFD : pic_data = 24'h956977;
          13'h1CFE : pic_data = 24'h956972;
          13'h1CFF : pic_data = 24'h956970;
          13'h1D00 : pic_data = 24'h95696e;
          13'h1D01 : pic_data = 24'h906f6f;
          13'h1D02 : pic_data = 24'h90706f;
          13'h1D03 : pic_data = 24'h90726f;
          13'h1D04 : pic_data = 24'h90756f;
          13'h1D05 : pic_data = 24'h90776f;
          13'h1D06 : pic_data = 24'h90796f;
          13'h1D07 : pic_data = 24'h90796f;
          13'h1D08 : pic_data = 24'h907b6f;
          13'h1D09 : pic_data = 24'h90806f;
          13'h1D0A : pic_data = 24'h90806f;
          13'h1D0B : pic_data = 24'h90836f;
          13'h1D0C : pic_data = 24'h90836f;
          13'h1D0D : pic_data = 24'h90856f;
          13'h1D0E : pic_data = 24'h908a6f;
          13'h1D0F : pic_data = 24'h908a6f;
          13'h1D10 : pic_data = 24'h908c6f;
          13'h1D11 : pic_data = 24'h908e6f;
          13'h1D12 : pic_data = 24'h91906f;
          13'h1D13 : pic_data = 24'h8c906f;
          13'h1D14 : pic_data = 24'h8b906f;
          13'h1D15 : pic_data = 24'h8a906f;
          13'h1D16 : pic_data = 24'h85906f;
          13'h1D17 : pic_data = 24'h86906f;
          13'h1D18 : pic_data = 24'h82906f;
          13'h1D19 : pic_data = 24'h82906f;
          13'h1D1A : pic_data = 24'h80906f;
          13'h1D1B : pic_data = 24'h7c906f;
          13'h1D1C : pic_data = 24'h7c906f;
          13'h1D1D : pic_data = 24'h78906f;
          13'h1D1E : pic_data = 24'h78906f;
          13'h1D1F : pic_data = 24'h75906f;
          13'h1D20 : pic_data = 24'h71906f;
          13'h1D21 : pic_data = 24'h72906f;
          13'h1D22 : pic_data = 24'h70906f;
          13'h1D23 : pic_data = 24'h6f9070;
          13'h1D24 : pic_data = 24'h6f9072;
          13'h1D25 : pic_data = 24'h6f9074;
          13'h1D26 : pic_data = 24'h6f9076;
          13'h1D27 : pic_data = 24'h6f9079;
          13'h1D28 : pic_data = 24'h6f907a;
          13'h1D29 : pic_data = 24'h6f907b;
          13'h1D2A : pic_data = 24'h6f907f;
          13'h1D2B : pic_data = 24'h6f9081;
          13'h1D2C : pic_data = 24'h6f9083;
          13'h1D2D : pic_data = 24'h6f9083;
          13'h1D2E : pic_data = 24'h6f9085;
          13'h1D2F : pic_data = 24'h6f9088;
          13'h1D30 : pic_data = 24'h6f908a;
          13'h1D31 : pic_data = 24'h6f908c;
          13'h1D32 : pic_data = 24'h6f908d;
          13'h1D33 : pic_data = 24'h6f9090;
          13'h1D34 : pic_data = 24'h6f8d90;
          13'h1D35 : pic_data = 24'h6f8b90;
          13'h1D36 : pic_data = 24'h6f8990;
          13'h1D37 : pic_data = 24'h6f8690;
          13'h1D38 : pic_data = 24'h6f8590;
          13'h1D39 : pic_data = 24'h6f8390;
          13'h1D3A : pic_data = 24'h6f8190;
          13'h1D3B : pic_data = 24'h6f8090;
          13'h1D3C : pic_data = 24'h6f7c90;
          13'h1D3D : pic_data = 24'h6f7c90;
          13'h1D3E : pic_data = 24'h6f7a90;
          13'h1D3F : pic_data = 24'h6f7890;
          13'h1D40 : pic_data = 24'h6f7590;
          13'h1D41 : pic_data = 24'h6f7390;
          13'h1D42 : pic_data = 24'h6f7290;
          13'h1D43 : pic_data = 24'h6f7090;
          13'h1D44 : pic_data = 24'h6f6f90;
          13'h1D45 : pic_data = 24'h726f90;
          13'h1D46 : pic_data = 24'h746f90;
          13'h1D47 : pic_data = 24'h766f90;
          13'h1D48 : pic_data = 24'h796f90;
          13'h1D49 : pic_data = 24'h786f90;
          13'h1D4A : pic_data = 24'h7c6f90;
          13'h1D4B : pic_data = 24'h7e6f90;
          13'h1D4C : pic_data = 24'h7f6f90;
          13'h1D4D : pic_data = 24'h836f90;
          13'h1D4E : pic_data = 24'h826f90;
          13'h1D4F : pic_data = 24'h856f90;
          13'h1D50 : pic_data = 24'h876f90;
          13'h1D51 : pic_data = 24'h896f90;
          13'h1D52 : pic_data = 24'h8c6f90;
          13'h1D53 : pic_data = 24'h8c6f90;
          13'h1D54 : pic_data = 24'h916f90;
          13'h1D55 : pic_data = 24'h906f8e;
          13'h1D56 : pic_data = 24'h906f8c;
          13'h1D57 : pic_data = 24'h906f89;
          13'h1D58 : pic_data = 24'h906f87;
          13'h1D59 : pic_data = 24'h906f85;
          13'h1D5A : pic_data = 24'h906f83;
          13'h1D5B : pic_data = 24'h906f83;
          13'h1D5C : pic_data = 24'h906f7f;
          13'h1D5D : pic_data = 24'h906f7e;
          13'h1D5E : pic_data = 24'h906f7c;
          13'h1D5F : pic_data = 24'h906f79;
          13'h1D60 : pic_data = 24'h906f79;
          13'h1D61 : pic_data = 24'h906f74;
          13'h1D62 : pic_data = 24'h906f73;
          13'h1D63 : pic_data = 24'h906f72;
          13'h1D64 : pic_data = 24'h916e6e;
          13'h1D65 : pic_data = 24'h916f6e;
          13'h1D66 : pic_data = 24'h91716e;
          13'h1D67 : pic_data = 24'h91746e;
          13'h1D68 : pic_data = 24'h91766e;
          13'h1D69 : pic_data = 24'h91796e;
          13'h1D6A : pic_data = 24'h91796e;
          13'h1D6B : pic_data = 24'h917b6e;
          13'h1D6C : pic_data = 24'h91806e;
          13'h1D6D : pic_data = 24'h91806e;
          13'h1D6E : pic_data = 24'h91836e;
          13'h1D6F : pic_data = 24'h91836e;
          13'h1D70 : pic_data = 24'h91856e;
          13'h1D71 : pic_data = 24'h918a6e;
          13'h1D72 : pic_data = 24'h918b6e;
          13'h1D73 : pic_data = 24'h918d6e;
          13'h1D74 : pic_data = 24'h918f6e;
          13'h1D75 : pic_data = 24'h91916e;
          13'h1D76 : pic_data = 24'h8c916e;
          13'h1D77 : pic_data = 24'h8c916e;
          13'h1D78 : pic_data = 24'h8a916e;
          13'h1D79 : pic_data = 24'h85916e;
          13'h1D7A : pic_data = 24'h86916e;
          13'h1D7B : pic_data = 24'h82916e;
          13'h1D7C : pic_data = 24'h82916e;
          13'h1D7D : pic_data = 24'h80916e;
          13'h1D7E : pic_data = 24'h7c916e;
          13'h1D7F : pic_data = 24'h7c916e;
          13'h1D80 : pic_data = 24'h78916e;
          13'h1D81 : pic_data = 24'h78916e;
          13'h1D82 : pic_data = 24'h74916e;
          13'h1D83 : pic_data = 24'h71916e;
          13'h1D84 : pic_data = 24'h72916e;
          13'h1D85 : pic_data = 24'h6f916e;
          13'h1D86 : pic_data = 24'h6e916f;
          13'h1D87 : pic_data = 24'h6e9171;
          13'h1D88 : pic_data = 24'h6e9173;
          13'h1D89 : pic_data = 24'h6e9175;
          13'h1D8A : pic_data = 24'h6e9179;
          13'h1D8B : pic_data = 24'h6e9179;
          13'h1D8C : pic_data = 24'h6e917b;
          13'h1D8D : pic_data = 24'h6e917f;
          13'h1D8E : pic_data = 24'h6e9181;
          13'h1D8F : pic_data = 24'h6e9183;
          13'h1D90 : pic_data = 24'h6e9183;
          13'h1D91 : pic_data = 24'h6e9185;
          13'h1D92 : pic_data = 24'h6e9189;
          13'h1D93 : pic_data = 24'h6e918b;
          13'h1D94 : pic_data = 24'h6e918d;
          13'h1D95 : pic_data = 24'h6e918e;
          13'h1D96 : pic_data = 24'h6e9191;
          13'h1D97 : pic_data = 24'h6e8e91;
          13'h1D98 : pic_data = 24'h6e8c91;
          13'h1D99 : pic_data = 24'h6e8a91;
          13'h1D9A : pic_data = 24'h6e8691;
          13'h1D9B : pic_data = 24'h6e8691;
          13'h1D9C : pic_data = 24'h6e8491;
          13'h1D9D : pic_data = 24'h6e8291;
          13'h1D9E : pic_data = 24'h6e8091;
          13'h1D9F : pic_data = 24'h6e7c91;
          13'h1DA0 : pic_data = 24'h6e7c91;
          13'h1DA1 : pic_data = 24'h6e7991;
          13'h1DA2 : pic_data = 24'h6e7791;
          13'h1DA3 : pic_data = 24'h6e7491;
          13'h1DA4 : pic_data = 24'h6e7291;
          13'h1DA5 : pic_data = 24'h6e7191;
          13'h1DA6 : pic_data = 24'h6e6f91;
          13'h1DA7 : pic_data = 24'h6e6e91;
          13'h1DA8 : pic_data = 24'h716e91;
          13'h1DA9 : pic_data = 24'h736e91;
          13'h1DAA : pic_data = 24'h756e91;
          13'h1DAB : pic_data = 24'h796e91;
          13'h1DAC : pic_data = 24'h786e91;
          13'h1DAD : pic_data = 24'h7c6e91;
          13'h1DAE : pic_data = 24'h7d6e91;
          13'h1DAF : pic_data = 24'h7f6e91;
          13'h1DB0 : pic_data = 24'h836e91;
          13'h1DB1 : pic_data = 24'h826e91;
          13'h1DB2 : pic_data = 24'h866e91;
          13'h1DB3 : pic_data = 24'h886e91;
          13'h1DB4 : pic_data = 24'h8a6e91;
          13'h1DB5 : pic_data = 24'h8d6e91;
          13'h1DB6 : pic_data = 24'h8c6e91;
          13'h1DB7 : pic_data = 24'h916e91;
          13'h1DB8 : pic_data = 24'h916e8f;
          13'h1DB9 : pic_data = 24'h916e8d;
          13'h1DBA : pic_data = 24'h916e8a;
          13'h1DBB : pic_data = 24'h916e88;
          13'h1DBC : pic_data = 24'h916e86;
          13'h1DBD : pic_data = 24'h916e83;
          13'h1DBE : pic_data = 24'h916e83;
          13'h1DBF : pic_data = 24'h916e7f;
          13'h1DC0 : pic_data = 24'h916e7e;
          13'h1DC1 : pic_data = 24'h916e7b;
          13'h1DC2 : pic_data = 24'h916e79;
          13'h1DC3 : pic_data = 24'h916e79;
          13'h1DC4 : pic_data = 24'h916e74;
          13'h1DC5 : pic_data = 24'h916e72;
          13'h1DC6 : pic_data = 24'h916e71;
          13'h1DC7 : pic_data = 24'h8e7071;
          13'h1DC8 : pic_data = 24'h8e7271;
          13'h1DC9 : pic_data = 24'h8e7371;
          13'h1DCA : pic_data = 24'h8e7671;
          13'h1DCB : pic_data = 24'h8e7871;
          13'h1DCC : pic_data = 24'h8e7971;
          13'h1DCD : pic_data = 24'h8e7a71;
          13'h1DCE : pic_data = 24'h8e7c71;
          13'h1DCF : pic_data = 24'h8e8071;
          13'h1DD0 : pic_data = 24'h8e8071;
          13'h1DD1 : pic_data = 24'h8e8271;
          13'h1DD2 : pic_data = 24'h8e8371;
          13'h1DD3 : pic_data = 24'h8e8571;
          13'h1DD4 : pic_data = 24'h8e8871;
          13'h1DD5 : pic_data = 24'h8e8971;
          13'h1DD6 : pic_data = 24'h8e8b71;
          13'h1DD7 : pic_data = 24'h8e8c71;
          13'h1DD8 : pic_data = 24'h8e8e71;
          13'h1DD9 : pic_data = 24'h8b8e71;
          13'h1DDA : pic_data = 24'h8a8e71;
          13'h1DDB : pic_data = 24'h888e71;
          13'h1DDC : pic_data = 24'h858e71;
          13'h1DDD : pic_data = 24'h858e71;
          13'h1DDE : pic_data = 24'h828e71;
          13'h1DDF : pic_data = 24'h818e71;
          13'h1DE0 : pic_data = 24'h808e71;
          13'h1DE1 : pic_data = 24'h7c8e71;
          13'h1DE2 : pic_data = 24'h7c8e71;
          13'h1DE3 : pic_data = 24'h798e71;
          13'h1DE4 : pic_data = 24'h788e71;
          13'h1DE5 : pic_data = 24'h768e71;
          13'h1DE6 : pic_data = 24'h738e71;
          13'h1DE7 : pic_data = 24'h738e71;
          13'h1DE8 : pic_data = 24'h718e70;
          13'h1DE9 : pic_data = 24'h718e72;
          13'h1DEA : pic_data = 24'h718e73;
          13'h1DEB : pic_data = 24'h718e75;
          13'h1DEC : pic_data = 24'h718e77;
          13'h1DED : pic_data = 24'h718e79;
          13'h1DEE : pic_data = 24'h718e7a;
          13'h1DEF : pic_data = 24'h718e7c;
          13'h1DF0 : pic_data = 24'h718e7f;
          13'h1DF1 : pic_data = 24'h718e81;
          13'h1DF2 : pic_data = 24'h718e82;
          13'h1DF3 : pic_data = 24'h718e83;
          13'h1DF4 : pic_data = 24'h718e85;
          13'h1DF5 : pic_data = 24'h718e88;
          13'h1DF6 : pic_data = 24'h718e89;
          13'h1DF7 : pic_data = 24'h718e8b;
          13'h1DF8 : pic_data = 24'h718e8b;
          13'h1DF9 : pic_data = 24'h718e8e;
          13'h1DFA : pic_data = 24'h718c8e;
          13'h1DFB : pic_data = 24'h718a8e;
          13'h1DFC : pic_data = 24'h71888e;
          13'h1DFD : pic_data = 24'h71868e;
          13'h1DFE : pic_data = 24'h71858e;
          13'h1DFF : pic_data = 24'h71838e;
          13'h1E00 : pic_data = 24'h71828e;
          13'h1E01 : pic_data = 24'h71808e;
          13'h1E02 : pic_data = 24'h717d8e;
          13'h1E03 : pic_data = 24'h717c8e;
          13'h1E04 : pic_data = 24'h717a8e;
          13'h1E05 : pic_data = 24'h71798e;
          13'h1E06 : pic_data = 24'h71768e;
          13'h1E07 : pic_data = 24'h71748e;
          13'h1E08 : pic_data = 24'h71738e;
          13'h1E09 : pic_data = 24'h71728e;
          13'h1E0A : pic_data = 24'h70708e;
          13'h1E0B : pic_data = 24'h73718e;
          13'h1E0C : pic_data = 24'h75718e;
          13'h1E0D : pic_data = 24'h76718e;
          13'h1E0E : pic_data = 24'h79718e;
          13'h1E0F : pic_data = 24'h79718e;
          13'h1E10 : pic_data = 24'h7c718e;
          13'h1E11 : pic_data = 24'h7e718e;
          13'h1E12 : pic_data = 24'h7f718e;
          13'h1E13 : pic_data = 24'h82718e;
          13'h1E14 : pic_data = 24'h82718e;
          13'h1E15 : pic_data = 24'h85718e;
          13'h1E16 : pic_data = 24'h86718e;
          13'h1E17 : pic_data = 24'h88718e;
          13'h1E18 : pic_data = 24'h8b718e;
          13'h1E19 : pic_data = 24'h8b718e;
          13'h1E1A : pic_data = 24'h8e718e;
          13'h1E1B : pic_data = 24'h8e718c;
          13'h1E1C : pic_data = 24'h8e718b;
          13'h1E1D : pic_data = 24'h8e7188;
          13'h1E1E : pic_data = 24'h8e7186;
          13'h1E1F : pic_data = 24'h8e7185;
          13'h1E20 : pic_data = 24'h8e7183;
          13'h1E21 : pic_data = 24'h8e7182;
          13'h1E22 : pic_data = 24'h8e717f;
          13'h1E23 : pic_data = 24'h8e717d;
          13'h1E24 : pic_data = 24'h8e717c;
          13'h1E25 : pic_data = 24'h8e717a;
          13'h1E26 : pic_data = 24'h8e7179;
          13'h1E27 : pic_data = 24'h8e7176;
          13'h1E28 : pic_data = 24'h8e7174;
          13'h1E29 : pic_data = 24'h8e7173;
          13'h1E2A : pic_data = 24'h8b7373;
          13'h1E2B : pic_data = 24'h8b7473;
          13'h1E2C : pic_data = 24'h8b7473;
          13'h1E2D : pic_data = 24'h8b7873;
          13'h1E2E : pic_data = 24'h8b7973;
          13'h1E2F : pic_data = 24'h8b7a73;
          13'h1E30 : pic_data = 24'h8b7a73;
          13'h1E31 : pic_data = 24'h8b7c73;
          13'h1E32 : pic_data = 24'h8b8073;
          13'h1E33 : pic_data = 24'h8b8173;
          13'h1E34 : pic_data = 24'h8b8173;
          13'h1E35 : pic_data = 24'h8b8273;
          13'h1E36 : pic_data = 24'h8b8473;
          13'h1E37 : pic_data = 24'h8b8673;
          13'h1E38 : pic_data = 24'h8b8773;
          13'h1E39 : pic_data = 24'h8b8973;
          13'h1E3A : pic_data = 24'h8b8a73;
          13'h1E3B : pic_data = 24'h8b8b73;
          13'h1E3C : pic_data = 24'h898b73;
          13'h1E3D : pic_data = 24'h888b73;
          13'h1E3E : pic_data = 24'h868b73;
          13'h1E3F : pic_data = 24'h848b73;
          13'h1E40 : pic_data = 24'h858b73;
          13'h1E41 : pic_data = 24'h818b73;
          13'h1E42 : pic_data = 24'h808b73;
          13'h1E43 : pic_data = 24'h808b73;
          13'h1E44 : pic_data = 24'h7c8b73;
          13'h1E45 : pic_data = 24'h7d8b73;
          13'h1E46 : pic_data = 24'h798b73;
          13'h1E47 : pic_data = 24'h798b73;
          13'h1E48 : pic_data = 24'h788b73;
          13'h1E49 : pic_data = 24'h748b73;
          13'h1E4A : pic_data = 24'h758b73;
          13'h1E4B : pic_data = 24'h728b73;
          13'h1E4C : pic_data = 24'h738b74;
          13'h1E4D : pic_data = 24'h738b75;
          13'h1E4E : pic_data = 24'h738b77;
          13'h1E4F : pic_data = 24'h738b79;
          13'h1E50 : pic_data = 24'h738b7a;
          13'h1E51 : pic_data = 24'h738b7a;
          13'h1E52 : pic_data = 24'h738b7d;
          13'h1E53 : pic_data = 24'h738b7f;
          13'h1E54 : pic_data = 24'h738b81;
          13'h1E55 : pic_data = 24'h738b81;
          13'h1E56 : pic_data = 24'h738b82;
          13'h1E57 : pic_data = 24'h738b84;
          13'h1E58 : pic_data = 24'h738b87;
          13'h1E59 : pic_data = 24'h738b87;
          13'h1E5A : pic_data = 24'h738b8a;
          13'h1E5B : pic_data = 24'h738b89;
          13'h1E5C : pic_data = 24'h738b8b;
          13'h1E5D : pic_data = 24'h738a8b;
          13'h1E5E : pic_data = 24'h73888b;
          13'h1E5F : pic_data = 24'h73868b;
          13'h1E60 : pic_data = 24'h73858b;
          13'h1E61 : pic_data = 24'h73858b;
          13'h1E62 : pic_data = 24'h73828b;
          13'h1E63 : pic_data = 24'h73828b;
          13'h1E64 : pic_data = 24'h73808b;
          13'h1E65 : pic_data = 24'h737d8b;
          13'h1E66 : pic_data = 24'h737d8b;
          13'h1E67 : pic_data = 24'h737a8b;
          13'h1E68 : pic_data = 24'h737a8b;
          13'h1E69 : pic_data = 24'h73788b;
          13'h1E6A : pic_data = 24'h73768b;
          13'h1E6B : pic_data = 24'h73758b;
          13'h1E6C : pic_data = 24'h73748b;
          13'h1E6D : pic_data = 24'h72738b;
          13'h1E6E : pic_data = 24'h75738b;
          13'h1E6F : pic_data = 24'h77738b;
          13'h1E70 : pic_data = 24'h77738b;
          13'h1E71 : pic_data = 24'h7a738b;
          13'h1E72 : pic_data = 24'h79738b;
          13'h1E73 : pic_data = 24'h7d738b;
          13'h1E74 : pic_data = 24'h7f738b;
          13'h1E75 : pic_data = 24'h7f738b;
          13'h1E76 : pic_data = 24'h82738b;
          13'h1E77 : pic_data = 24'h81738b;
          13'h1E78 : pic_data = 24'h85738b;
          13'h1E79 : pic_data = 24'h85738b;
          13'h1E7A : pic_data = 24'h86738b;
          13'h1E7B : pic_data = 24'h8a738b;
          13'h1E7C : pic_data = 24'h89738b;
          13'h1E7D : pic_data = 24'h8b738b;
          13'h1E7E : pic_data = 24'h8b738a;
          13'h1E7F : pic_data = 24'h8b738a;
          13'h1E80 : pic_data = 24'h8b7386;
          13'h1E81 : pic_data = 24'h8b7385;
          13'h1E82 : pic_data = 24'h8b7385;
          13'h1E83 : pic_data = 24'h8b7382;
          13'h1E84 : pic_data = 24'h8b7382;
          13'h1E85 : pic_data = 24'h8b7380;
          13'h1E86 : pic_data = 24'h8b737d;
          13'h1E87 : pic_data = 24'h8b737d;
          13'h1E88 : pic_data = 24'h8b737a;
          13'h1E89 : pic_data = 24'h8b737a;
          13'h1E8A : pic_data = 24'h8b7378;
          13'h1E8B : pic_data = 24'h8b7376;
          13'h1E8C : pic_data = 24'h8b7375;
          13'h1E8D : pic_data = 24'h8c7273;
          13'h1E8E : pic_data = 24'h8c7473;
          13'h1E8F : pic_data = 24'h8c7473;
          13'h1E90 : pic_data = 24'h8c7873;
          13'h1E91 : pic_data = 24'h8c7973;
          13'h1E92 : pic_data = 24'h8c7a73;
          13'h1E93 : pic_data = 24'h8c7a73;
          13'h1E94 : pic_data = 24'h8c7c73;
          13'h1E95 : pic_data = 24'h8c8073;
          13'h1E96 : pic_data = 24'h8c8173;
          13'h1E97 : pic_data = 24'h8c8273;
          13'h1E98 : pic_data = 24'h8c8273;
          13'h1E99 : pic_data = 24'h8c8573;
          13'h1E9A : pic_data = 24'h8c8773;
          13'h1E9B : pic_data = 24'h8c8773;
          13'h1E9C : pic_data = 24'h8c8a73;
          13'h1E9D : pic_data = 24'h8c8b73;
          13'h1E9E : pic_data = 24'h8c8c73;
          13'h1E9F : pic_data = 24'h898c73;
          13'h1EA0 : pic_data = 24'h898c73;
          13'h1EA1 : pic_data = 24'h878c73;
          13'h1EA2 : pic_data = 24'h848c73;
          13'h1EA3 : pic_data = 24'h858c73;
          13'h1EA4 : pic_data = 24'h818c73;
          13'h1EA5 : pic_data = 24'h818c73;
          13'h1EA6 : pic_data = 24'h808c73;
          13'h1EA7 : pic_data = 24'h7c8c73;
          13'h1EA8 : pic_data = 24'h7d8c73;
          13'h1EA9 : pic_data = 24'h798c73;
          13'h1EAA : pic_data = 24'h798c73;
          13'h1EAB : pic_data = 24'h788c73;
          13'h1EAC : pic_data = 24'h748c73;
          13'h1EAD : pic_data = 24'h758c73;
          13'h1EAE : pic_data = 24'h728c72;
          13'h1EAF : pic_data = 24'h738c74;
          13'h1EB0 : pic_data = 24'h738c74;
          13'h1EB1 : pic_data = 24'h738c77;
          13'h1EB2 : pic_data = 24'h738c79;
          13'h1EB3 : pic_data = 24'h738c7a;
          13'h1EB4 : pic_data = 24'h738c7a;
          13'h1EB5 : pic_data = 24'h738c7d;
          13'h1EB6 : pic_data = 24'h738c7f;
          13'h1EB7 : pic_data = 24'h738c81;
          13'h1EB8 : pic_data = 24'h738c82;
          13'h1EB9 : pic_data = 24'h738c82;
          13'h1EBA : pic_data = 24'h738c85;
          13'h1EBB : pic_data = 24'h738c87;
          13'h1EBC : pic_data = 24'h738c87;
          13'h1EBD : pic_data = 24'h738c8a;
          13'h1EBE : pic_data = 24'h738c89;
          13'h1EBF : pic_data = 24'h738c8c;
          13'h1EC0 : pic_data = 24'h738b8c;
          13'h1EC1 : pic_data = 24'h73898c;
          13'h1EC2 : pic_data = 24'h73868c;
          13'h1EC3 : pic_data = 24'h73868c;
          13'h1EC4 : pic_data = 24'h73858c;
          13'h1EC5 : pic_data = 24'h73828c;
          13'h1EC6 : pic_data = 24'h73828c;
          13'h1EC7 : pic_data = 24'h73808c;
          13'h1EC8 : pic_data = 24'h737d8c;
          13'h1EC9 : pic_data = 24'h737d8c;
          13'h1ECA : pic_data = 24'h737a8c;
          13'h1ECB : pic_data = 24'h737a8c;
          13'h1ECC : pic_data = 24'h73788c;
          13'h1ECD : pic_data = 24'h73758c;
          13'h1ECE : pic_data = 24'h73758c;
          13'h1ECF : pic_data = 24'h73748c;
          13'h1ED0 : pic_data = 24'h72728c;
          13'h1ED1 : pic_data = 24'h75738c;
          13'h1ED2 : pic_data = 24'h77738c;
          13'h1ED3 : pic_data = 24'h77738c;
          13'h1ED4 : pic_data = 24'h7a738c;
          13'h1ED5 : pic_data = 24'h79738c;
          13'h1ED6 : pic_data = 24'h7d738c;
          13'h1ED7 : pic_data = 24'h7f738c;
          13'h1ED8 : pic_data = 24'h7f738c;
          13'h1ED9 : pic_data = 24'h82738c;
          13'h1EDA : pic_data = 24'h81738c;
          13'h1EDB : pic_data = 24'h85738c;
          13'h1EDC : pic_data = 24'h86738c;
          13'h1EDD : pic_data = 24'h86738c;
          13'h1EDE : pic_data = 24'h8a738c;
          13'h1EDF : pic_data = 24'h89738c;
          13'h1EE0 : pic_data = 24'h8c738c;
          13'h1EE1 : pic_data = 24'h8c738b;
          13'h1EE2 : pic_data = 24'h8c738a;
          13'h1EE3 : pic_data = 24'h8c7386;
          13'h1EE4 : pic_data = 24'h8c7386;
          13'h1EE5 : pic_data = 24'h8c7385;
          13'h1EE6 : pic_data = 24'h8c7382;
          13'h1EE7 : pic_data = 24'h8c7382;
          13'h1EE8 : pic_data = 24'h8c7380;
          13'h1EE9 : pic_data = 24'h8c737d;
          13'h1EEA : pic_data = 24'h8c737d;
          13'h1EEB : pic_data = 24'h8c737a;
          13'h1EEC : pic_data = 24'h8c737a;
          13'h1EED : pic_data = 24'h8c7378;
          13'h1EEE : pic_data = 24'h8c7375;
          default  : pic_data = 24'h8c7374;
      endcase
  end
`elsif TEST_PAT2
  always @(*) begin
      pic_data = hcnt ^ vcnt;
  end
`elsif TEST_PAT3
  always @(*) begin
      case (hcnt[8:7] + vcnt[8:7])
          3'h0   : pic_data = 24'hFF0000;
          3'h1   : pic_data = 24'h00FF00;
          3'h2   : pic_data = 24'h0000FF;
          3'h3   : pic_data = 24'h808000;
          3'h4   : pic_data = 24'h008080;
          3'h5   : pic_data = 24'h800080;
          default: pic_data = 24'hFFFFFF;
      endcase
  end
`endif

  assign pic_hsync = (hcnt == 0) | ((hcnt > 0) & (hcnt <= (HSTART - 10)));
  assign pic_vsync = (vcnt == 0) | ((vcnt > 0) & (vcnt <= (VSTART - 10)));

endmodule
